module PreDecode_top;

  wire [15:0] io_in_bits_data_0;
  wire [15:0] io_in_bits_data_1;
  wire [15:0] io_in_bits_data_2;
  wire [15:0] io_in_bits_data_3;
  wire [15:0] io_in_bits_data_4;
  wire [15:0] io_in_bits_data_5;
  wire [15:0] io_in_bits_data_6;
  wire [15:0] io_in_bits_data_7;
  wire [15:0] io_in_bits_data_8;
  wire [15:0] io_in_bits_data_9;
  wire [15:0] io_in_bits_data_10;
  wire [15:0] io_in_bits_data_11;
  wire [15:0] io_in_bits_data_12;
  wire [15:0] io_in_bits_data_13;
  wire [15:0] io_in_bits_data_14;
  wire [15:0] io_in_bits_data_15;
  wire [15:0] io_in_bits_data_16;
  wire  io_out_pd_0_isRVC;
  wire  io_out_pd_1_valid;
  wire  io_out_pd_1_isRVC;
  wire  io_out_pd_2_valid;
  wire  io_out_pd_2_isRVC;
  wire  io_out_pd_3_valid;
  wire  io_out_pd_3_isRVC;
  wire  io_out_pd_4_valid;
  wire  io_out_pd_4_isRVC;
  wire  io_out_pd_5_valid;
  wire  io_out_pd_5_isRVC;
  wire  io_out_pd_6_valid;
  wire  io_out_pd_6_isRVC;
  wire  io_out_pd_7_valid;
  wire  io_out_pd_7_isRVC;
  wire  io_out_pd_8_valid;
  wire  io_out_pd_8_isRVC;
  wire  io_out_pd_9_valid;
  wire  io_out_pd_9_isRVC;
  wire  io_out_pd_10_valid;
  wire  io_out_pd_10_isRVC;
  wire  io_out_pd_11_valid;
  wire  io_out_pd_11_isRVC;
  wire  io_out_pd_12_valid;
  wire  io_out_pd_12_isRVC;
  wire  io_out_pd_13_valid;
  wire  io_out_pd_13_isRVC;
  wire  io_out_pd_14_valid;
  wire  io_out_pd_14_isRVC;
  wire  io_out_pd_15_valid;
  wire  io_out_pd_15_isRVC;
  wire  io_out_hasHalfValid_2;
  wire  io_out_hasHalfValid_3;
  wire  io_out_hasHalfValid_4;
  wire  io_out_hasHalfValid_5;
  wire  io_out_hasHalfValid_6;
  wire  io_out_hasHalfValid_7;
  wire  io_out_hasHalfValid_8;
  wire  io_out_hasHalfValid_9;
  wire  io_out_hasHalfValid_10;
  wire  io_out_hasHalfValid_11;
  wire  io_out_hasHalfValid_12;
  wire  io_out_hasHalfValid_13;
  wire  io_out_hasHalfValid_14;
  wire  io_out_hasHalfValid_15;
  wire [31:0] io_out_instr_0;
  wire [31:0] io_out_instr_1;
  wire [31:0] io_out_instr_2;
  wire [31:0] io_out_instr_3;
  wire [31:0] io_out_instr_4;
  wire [31:0] io_out_instr_5;
  wire [31:0] io_out_instr_6;
  wire [31:0] io_out_instr_7;
  wire [31:0] io_out_instr_8;
  wire [31:0] io_out_instr_9;
  wire [31:0] io_out_instr_10;
  wire [31:0] io_out_instr_11;
  wire [31:0] io_out_instr_12;
  wire [31:0] io_out_instr_13;
  wire [31:0] io_out_instr_14;
  wire [31:0] io_out_instr_15;
  wire [63:0] io_out_jumpOffset_0;
  wire [63:0] io_out_jumpOffset_1;
  wire [63:0] io_out_jumpOffset_2;
  wire [63:0] io_out_jumpOffset_3;
  wire [63:0] io_out_jumpOffset_4;
  wire [63:0] io_out_jumpOffset_5;
  wire [63:0] io_out_jumpOffset_6;
  wire [63:0] io_out_jumpOffset_7;
  wire [63:0] io_out_jumpOffset_8;
  wire [63:0] io_out_jumpOffset_9;
  wire [63:0] io_out_jumpOffset_10;
  wire [63:0] io_out_jumpOffset_11;
  wire [63:0] io_out_jumpOffset_12;
  wire [63:0] io_out_jumpOffset_13;
  wire [63:0] io_out_jumpOffset_14;
  wire [63:0] io_out_jumpOffset_15;


 PreDecode PreDecode(
    .io_in_bits_data_0(io_in_bits_data_0),
    .io_in_bits_data_1(io_in_bits_data_1),
    .io_in_bits_data_2(io_in_bits_data_2),
    .io_in_bits_data_3(io_in_bits_data_3),
    .io_in_bits_data_4(io_in_bits_data_4),
    .io_in_bits_data_5(io_in_bits_data_5),
    .io_in_bits_data_6(io_in_bits_data_6),
    .io_in_bits_data_7(io_in_bits_data_7),
    .io_in_bits_data_8(io_in_bits_data_8),
    .io_in_bits_data_9(io_in_bits_data_9),
    .io_in_bits_data_10(io_in_bits_data_10),
    .io_in_bits_data_11(io_in_bits_data_11),
    .io_in_bits_data_12(io_in_bits_data_12),
    .io_in_bits_data_13(io_in_bits_data_13),
    .io_in_bits_data_14(io_in_bits_data_14),
    .io_in_bits_data_15(io_in_bits_data_15),
    .io_in_bits_data_16(io_in_bits_data_16),
    .io_out_pd_0_isRVC(io_out_pd_0_isRVC),
    .io_out_pd_1_valid(io_out_pd_1_valid),
    .io_out_pd_1_isRVC(io_out_pd_1_isRVC),
    .io_out_pd_2_valid(io_out_pd_2_valid),
    .io_out_pd_2_isRVC(io_out_pd_2_isRVC),
    .io_out_pd_3_valid(io_out_pd_3_valid),
    .io_out_pd_3_isRVC(io_out_pd_3_isRVC),
    .io_out_pd_4_valid(io_out_pd_4_valid),
    .io_out_pd_4_isRVC(io_out_pd_4_isRVC),
    .io_out_pd_5_valid(io_out_pd_5_valid),
    .io_out_pd_5_isRVC(io_out_pd_5_isRVC),
    .io_out_pd_6_valid(io_out_pd_6_valid),
    .io_out_pd_6_isRVC(io_out_pd_6_isRVC),
    .io_out_pd_7_valid(io_out_pd_7_valid),
    .io_out_pd_7_isRVC(io_out_pd_7_isRVC),
    .io_out_pd_8_valid(io_out_pd_8_valid),
    .io_out_pd_8_isRVC(io_out_pd_8_isRVC),
    .io_out_pd_9_valid(io_out_pd_9_valid),
    .io_out_pd_9_isRVC(io_out_pd_9_isRVC),
    .io_out_pd_10_valid(io_out_pd_10_valid),
    .io_out_pd_10_isRVC(io_out_pd_10_isRVC),
    .io_out_pd_11_valid(io_out_pd_11_valid),
    .io_out_pd_11_isRVC(io_out_pd_11_isRVC),
    .io_out_pd_12_valid(io_out_pd_12_valid),
    .io_out_pd_12_isRVC(io_out_pd_12_isRVC),
    .io_out_pd_13_valid(io_out_pd_13_valid),
    .io_out_pd_13_isRVC(io_out_pd_13_isRVC),
    .io_out_pd_14_valid(io_out_pd_14_valid),
    .io_out_pd_14_isRVC(io_out_pd_14_isRVC),
    .io_out_pd_15_valid(io_out_pd_15_valid),
    .io_out_pd_15_isRVC(io_out_pd_15_isRVC),
    .io_out_hasHalfValid_2(io_out_hasHalfValid_2),
    .io_out_hasHalfValid_3(io_out_hasHalfValid_3),
    .io_out_hasHalfValid_4(io_out_hasHalfValid_4),
    .io_out_hasHalfValid_5(io_out_hasHalfValid_5),
    .io_out_hasHalfValid_6(io_out_hasHalfValid_6),
    .io_out_hasHalfValid_7(io_out_hasHalfValid_7),
    .io_out_hasHalfValid_8(io_out_hasHalfValid_8),
    .io_out_hasHalfValid_9(io_out_hasHalfValid_9),
    .io_out_hasHalfValid_10(io_out_hasHalfValid_10),
    .io_out_hasHalfValid_11(io_out_hasHalfValid_11),
    .io_out_hasHalfValid_12(io_out_hasHalfValid_12),
    .io_out_hasHalfValid_13(io_out_hasHalfValid_13),
    .io_out_hasHalfValid_14(io_out_hasHalfValid_14),
    .io_out_hasHalfValid_15(io_out_hasHalfValid_15),
    .io_out_instr_0(io_out_instr_0),
    .io_out_instr_1(io_out_instr_1),
    .io_out_instr_2(io_out_instr_2),
    .io_out_instr_3(io_out_instr_3),
    .io_out_instr_4(io_out_instr_4),
    .io_out_instr_5(io_out_instr_5),
    .io_out_instr_6(io_out_instr_6),
    .io_out_instr_7(io_out_instr_7),
    .io_out_instr_8(io_out_instr_8),
    .io_out_instr_9(io_out_instr_9),
    .io_out_instr_10(io_out_instr_10),
    .io_out_instr_11(io_out_instr_11),
    .io_out_instr_12(io_out_instr_12),
    .io_out_instr_13(io_out_instr_13),
    .io_out_instr_14(io_out_instr_14),
    .io_out_instr_15(io_out_instr_15),
    .io_out_jumpOffset_0(io_out_jumpOffset_0),
    .io_out_jumpOffset_1(io_out_jumpOffset_1),
    .io_out_jumpOffset_2(io_out_jumpOffset_2),
    .io_out_jumpOffset_3(io_out_jumpOffset_3),
    .io_out_jumpOffset_4(io_out_jumpOffset_4),
    .io_out_jumpOffset_5(io_out_jumpOffset_5),
    .io_out_jumpOffset_6(io_out_jumpOffset_6),
    .io_out_jumpOffset_7(io_out_jumpOffset_7),
    .io_out_jumpOffset_8(io_out_jumpOffset_8),
    .io_out_jumpOffset_9(io_out_jumpOffset_9),
    .io_out_jumpOffset_10(io_out_jumpOffset_10),
    .io_out_jumpOffset_11(io_out_jumpOffset_11),
    .io_out_jumpOffset_12(io_out_jumpOffset_12),
    .io_out_jumpOffset_13(io_out_jumpOffset_13),
    .io_out_jumpOffset_14(io_out_jumpOffset_14),
    .io_out_jumpOffset_15(io_out_jumpOffset_15)
 );


endmodule

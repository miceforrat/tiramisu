module PredChecker_top;

  wire  clock;
  wire  io_in_ftqOffset_valid;
  wire [3:0] io_in_ftqOffset_bits;
  wire [63:0] io_in_jumpOffset_0;
  wire [63:0] io_in_jumpOffset_1;
  wire [63:0] io_in_jumpOffset_2;
  wire [63:0] io_in_jumpOffset_3;
  wire [63:0] io_in_jumpOffset_4;
  wire [63:0] io_in_jumpOffset_5;
  wire [63:0] io_in_jumpOffset_6;
  wire [63:0] io_in_jumpOffset_7;
  wire [63:0] io_in_jumpOffset_8;
  wire [63:0] io_in_jumpOffset_9;
  wire [63:0] io_in_jumpOffset_10;
  wire [63:0] io_in_jumpOffset_11;
  wire [63:0] io_in_jumpOffset_12;
  wire [63:0] io_in_jumpOffset_13;
  wire [63:0] io_in_jumpOffset_14;
  wire [63:0] io_in_jumpOffset_15;
  wire [49:0] io_in_target;
  wire  io_in_instrRange_0;
  wire  io_in_instrRange_1;
  wire  io_in_instrRange_2;
  wire  io_in_instrRange_3;
  wire  io_in_instrRange_4;
  wire  io_in_instrRange_5;
  wire  io_in_instrRange_6;
  wire  io_in_instrRange_7;
  wire  io_in_instrRange_8;
  wire  io_in_instrRange_9;
  wire  io_in_instrRange_10;
  wire  io_in_instrRange_11;
  wire  io_in_instrRange_12;
  wire  io_in_instrRange_13;
  wire  io_in_instrRange_14;
  wire  io_in_instrRange_15;
  wire  io_in_instrValid_0;
  wire  io_in_instrValid_1;
  wire  io_in_instrValid_2;
  wire  io_in_instrValid_3;
  wire  io_in_instrValid_4;
  wire  io_in_instrValid_5;
  wire  io_in_instrValid_6;
  wire  io_in_instrValid_7;
  wire  io_in_instrValid_8;
  wire  io_in_instrValid_9;
  wire  io_in_instrValid_10;
  wire  io_in_instrValid_11;
  wire  io_in_instrValid_12;
  wire  io_in_instrValid_13;
  wire  io_in_instrValid_14;
  wire  io_in_instrValid_15;
  wire  io_in_pds_0_isRVC;
  wire [1:0] io_in_pds_0_brType;
  wire  io_in_pds_0_isRet;
  wire  io_in_pds_1_isRVC;
  wire [1:0] io_in_pds_1_brType;
  wire  io_in_pds_1_isRet;
  wire  io_in_pds_2_isRVC;
  wire [1:0] io_in_pds_2_brType;
  wire  io_in_pds_2_isRet;
  wire  io_in_pds_3_isRVC;
  wire [1:0] io_in_pds_3_brType;
  wire  io_in_pds_3_isRet;
  wire  io_in_pds_4_isRVC;
  wire [1:0] io_in_pds_4_brType;
  wire  io_in_pds_4_isRet;
  wire  io_in_pds_5_isRVC;
  wire [1:0] io_in_pds_5_brType;
  wire  io_in_pds_5_isRet;
  wire  io_in_pds_6_isRVC;
  wire [1:0] io_in_pds_6_brType;
  wire  io_in_pds_6_isRet;
  wire  io_in_pds_7_isRVC;
  wire [1:0] io_in_pds_7_brType;
  wire  io_in_pds_7_isRet;
  wire  io_in_pds_8_isRVC;
  wire [1:0] io_in_pds_8_brType;
  wire  io_in_pds_8_isRet;
  wire  io_in_pds_9_isRVC;
  wire [1:0] io_in_pds_9_brType;
  wire  io_in_pds_9_isRet;
  wire  io_in_pds_10_isRVC;
  wire [1:0] io_in_pds_10_brType;
  wire  io_in_pds_10_isRet;
  wire  io_in_pds_11_isRVC;
  wire [1:0] io_in_pds_11_brType;
  wire  io_in_pds_11_isRet;
  wire  io_in_pds_12_isRVC;
  wire [1:0] io_in_pds_12_brType;
  wire  io_in_pds_12_isRet;
  wire  io_in_pds_13_isRVC;
  wire [1:0] io_in_pds_13_brType;
  wire  io_in_pds_13_isRet;
  wire  io_in_pds_14_isRVC;
  wire [1:0] io_in_pds_14_brType;
  wire  io_in_pds_14_isRet;
  wire  io_in_pds_15_isRVC;
  wire [1:0] io_in_pds_15_brType;
  wire  io_in_pds_15_isRet;
  wire [49:0] io_in_pc_0;
  wire [49:0] io_in_pc_1;
  wire [49:0] io_in_pc_2;
  wire [49:0] io_in_pc_3;
  wire [49:0] io_in_pc_4;
  wire [49:0] io_in_pc_5;
  wire [49:0] io_in_pc_6;
  wire [49:0] io_in_pc_7;
  wire [49:0] io_in_pc_8;
  wire [49:0] io_in_pc_9;
  wire [49:0] io_in_pc_10;
  wire [49:0] io_in_pc_11;
  wire [49:0] io_in_pc_12;
  wire [49:0] io_in_pc_13;
  wire [49:0] io_in_pc_14;
  wire [49:0] io_in_pc_15;
  wire  io_in_fire_in;
  wire  io_out_stage1Out_fixedRange_0;
  wire  io_out_stage1Out_fixedRange_1;
  wire  io_out_stage1Out_fixedRange_2;
  wire  io_out_stage1Out_fixedRange_3;
  wire  io_out_stage1Out_fixedRange_4;
  wire  io_out_stage1Out_fixedRange_5;
  wire  io_out_stage1Out_fixedRange_6;
  wire  io_out_stage1Out_fixedRange_7;
  wire  io_out_stage1Out_fixedRange_8;
  wire  io_out_stage1Out_fixedRange_9;
  wire  io_out_stage1Out_fixedRange_10;
  wire  io_out_stage1Out_fixedRange_11;
  wire  io_out_stage1Out_fixedRange_12;
  wire  io_out_stage1Out_fixedRange_13;
  wire  io_out_stage1Out_fixedRange_14;
  wire  io_out_stage1Out_fixedRange_15;
  wire  io_out_stage1Out_fixedTaken_0;
  wire  io_out_stage1Out_fixedTaken_1;
  wire  io_out_stage1Out_fixedTaken_2;
  wire  io_out_stage1Out_fixedTaken_3;
  wire  io_out_stage1Out_fixedTaken_4;
  wire  io_out_stage1Out_fixedTaken_5;
  wire  io_out_stage1Out_fixedTaken_6;
  wire  io_out_stage1Out_fixedTaken_7;
  wire  io_out_stage1Out_fixedTaken_8;
  wire  io_out_stage1Out_fixedTaken_9;
  wire  io_out_stage1Out_fixedTaken_10;
  wire  io_out_stage1Out_fixedTaken_11;
  wire  io_out_stage1Out_fixedTaken_12;
  wire  io_out_stage1Out_fixedTaken_13;
  wire  io_out_stage1Out_fixedTaken_14;
  wire  io_out_stage1Out_fixedTaken_15;
  wire [49:0] io_out_stage2Out_fixedTarget_0;
  wire [49:0] io_out_stage2Out_fixedTarget_1;
  wire [49:0] io_out_stage2Out_fixedTarget_2;
  wire [49:0] io_out_stage2Out_fixedTarget_3;
  wire [49:0] io_out_stage2Out_fixedTarget_4;
  wire [49:0] io_out_stage2Out_fixedTarget_5;
  wire [49:0] io_out_stage2Out_fixedTarget_6;
  wire [49:0] io_out_stage2Out_fixedTarget_7;
  wire [49:0] io_out_stage2Out_fixedTarget_8;
  wire [49:0] io_out_stage2Out_fixedTarget_9;
  wire [49:0] io_out_stage2Out_fixedTarget_10;
  wire [49:0] io_out_stage2Out_fixedTarget_11;
  wire [49:0] io_out_stage2Out_fixedTarget_12;
  wire [49:0] io_out_stage2Out_fixedTarget_13;
  wire [49:0] io_out_stage2Out_fixedTarget_14;
  wire [49:0] io_out_stage2Out_fixedTarget_15;
  wire [49:0] io_out_stage2Out_jalTarget_0;
  wire [49:0] io_out_stage2Out_jalTarget_1;
  wire [49:0] io_out_stage2Out_jalTarget_2;
  wire [49:0] io_out_stage2Out_jalTarget_3;
  wire [49:0] io_out_stage2Out_jalTarget_4;
  wire [49:0] io_out_stage2Out_jalTarget_5;
  wire [49:0] io_out_stage2Out_jalTarget_6;
  wire [49:0] io_out_stage2Out_jalTarget_7;
  wire [49:0] io_out_stage2Out_jalTarget_8;
  wire [49:0] io_out_stage2Out_jalTarget_9;
  wire [49:0] io_out_stage2Out_jalTarget_10;
  wire [49:0] io_out_stage2Out_jalTarget_11;
  wire [49:0] io_out_stage2Out_jalTarget_12;
  wire [49:0] io_out_stage2Out_jalTarget_13;
  wire [49:0] io_out_stage2Out_jalTarget_14;
  wire [49:0] io_out_stage2Out_jalTarget_15;
  wire  io_out_stage2Out_fixedMissPred_0;
  wire  io_out_stage2Out_fixedMissPred_1;
  wire  io_out_stage2Out_fixedMissPred_2;
  wire  io_out_stage2Out_fixedMissPred_3;
  wire  io_out_stage2Out_fixedMissPred_4;
  wire  io_out_stage2Out_fixedMissPred_5;
  wire  io_out_stage2Out_fixedMissPred_6;
  wire  io_out_stage2Out_fixedMissPred_7;
  wire  io_out_stage2Out_fixedMissPred_8;
  wire  io_out_stage2Out_fixedMissPred_9;
  wire  io_out_stage2Out_fixedMissPred_10;
  wire  io_out_stage2Out_fixedMissPred_11;
  wire  io_out_stage2Out_fixedMissPred_12;
  wire  io_out_stage2Out_fixedMissPred_13;
  wire  io_out_stage2Out_fixedMissPred_14;
  wire  io_out_stage2Out_fixedMissPred_15;


 PredChecker PredChecker(
    .clock(clock),
    .io_in_ftqOffset_valid(io_in_ftqOffset_valid),
    .io_in_ftqOffset_bits(io_in_ftqOffset_bits),
    .io_in_jumpOffset_0(io_in_jumpOffset_0),
    .io_in_jumpOffset_1(io_in_jumpOffset_1),
    .io_in_jumpOffset_2(io_in_jumpOffset_2),
    .io_in_jumpOffset_3(io_in_jumpOffset_3),
    .io_in_jumpOffset_4(io_in_jumpOffset_4),
    .io_in_jumpOffset_5(io_in_jumpOffset_5),
    .io_in_jumpOffset_6(io_in_jumpOffset_6),
    .io_in_jumpOffset_7(io_in_jumpOffset_7),
    .io_in_jumpOffset_8(io_in_jumpOffset_8),
    .io_in_jumpOffset_9(io_in_jumpOffset_9),
    .io_in_jumpOffset_10(io_in_jumpOffset_10),
    .io_in_jumpOffset_11(io_in_jumpOffset_11),
    .io_in_jumpOffset_12(io_in_jumpOffset_12),
    .io_in_jumpOffset_13(io_in_jumpOffset_13),
    .io_in_jumpOffset_14(io_in_jumpOffset_14),
    .io_in_jumpOffset_15(io_in_jumpOffset_15),
    .io_in_target(io_in_target),
    .io_in_instrRange_0(io_in_instrRange_0),
    .io_in_instrRange_1(io_in_instrRange_1),
    .io_in_instrRange_2(io_in_instrRange_2),
    .io_in_instrRange_3(io_in_instrRange_3),
    .io_in_instrRange_4(io_in_instrRange_4),
    .io_in_instrRange_5(io_in_instrRange_5),
    .io_in_instrRange_6(io_in_instrRange_6),
    .io_in_instrRange_7(io_in_instrRange_7),
    .io_in_instrRange_8(io_in_instrRange_8),
    .io_in_instrRange_9(io_in_instrRange_9),
    .io_in_instrRange_10(io_in_instrRange_10),
    .io_in_instrRange_11(io_in_instrRange_11),
    .io_in_instrRange_12(io_in_instrRange_12),
    .io_in_instrRange_13(io_in_instrRange_13),
    .io_in_instrRange_14(io_in_instrRange_14),
    .io_in_instrRange_15(io_in_instrRange_15),
    .io_in_instrValid_0(io_in_instrValid_0),
    .io_in_instrValid_1(io_in_instrValid_1),
    .io_in_instrValid_2(io_in_instrValid_2),
    .io_in_instrValid_3(io_in_instrValid_3),
    .io_in_instrValid_4(io_in_instrValid_4),
    .io_in_instrValid_5(io_in_instrValid_5),
    .io_in_instrValid_6(io_in_instrValid_6),
    .io_in_instrValid_7(io_in_instrValid_7),
    .io_in_instrValid_8(io_in_instrValid_8),
    .io_in_instrValid_9(io_in_instrValid_9),
    .io_in_instrValid_10(io_in_instrValid_10),
    .io_in_instrValid_11(io_in_instrValid_11),
    .io_in_instrValid_12(io_in_instrValid_12),
    .io_in_instrValid_13(io_in_instrValid_13),
    .io_in_instrValid_14(io_in_instrValid_14),
    .io_in_instrValid_15(io_in_instrValid_15),
    .io_in_pds_0_isRVC(io_in_pds_0_isRVC),
    .io_in_pds_0_brType(io_in_pds_0_brType),
    .io_in_pds_0_isRet(io_in_pds_0_isRet),
    .io_in_pds_1_isRVC(io_in_pds_1_isRVC),
    .io_in_pds_1_brType(io_in_pds_1_brType),
    .io_in_pds_1_isRet(io_in_pds_1_isRet),
    .io_in_pds_2_isRVC(io_in_pds_2_isRVC),
    .io_in_pds_2_brType(io_in_pds_2_brType),
    .io_in_pds_2_isRet(io_in_pds_2_isRet),
    .io_in_pds_3_isRVC(io_in_pds_3_isRVC),
    .io_in_pds_3_brType(io_in_pds_3_brType),
    .io_in_pds_3_isRet(io_in_pds_3_isRet),
    .io_in_pds_4_isRVC(io_in_pds_4_isRVC),
    .io_in_pds_4_brType(io_in_pds_4_brType),
    .io_in_pds_4_isRet(io_in_pds_4_isRet),
    .io_in_pds_5_isRVC(io_in_pds_5_isRVC),
    .io_in_pds_5_brType(io_in_pds_5_brType),
    .io_in_pds_5_isRet(io_in_pds_5_isRet),
    .io_in_pds_6_isRVC(io_in_pds_6_isRVC),
    .io_in_pds_6_brType(io_in_pds_6_brType),
    .io_in_pds_6_isRet(io_in_pds_6_isRet),
    .io_in_pds_7_isRVC(io_in_pds_7_isRVC),
    .io_in_pds_7_brType(io_in_pds_7_brType),
    .io_in_pds_7_isRet(io_in_pds_7_isRet),
    .io_in_pds_8_isRVC(io_in_pds_8_isRVC),
    .io_in_pds_8_brType(io_in_pds_8_brType),
    .io_in_pds_8_isRet(io_in_pds_8_isRet),
    .io_in_pds_9_isRVC(io_in_pds_9_isRVC),
    .io_in_pds_9_brType(io_in_pds_9_brType),
    .io_in_pds_9_isRet(io_in_pds_9_isRet),
    .io_in_pds_10_isRVC(io_in_pds_10_isRVC),
    .io_in_pds_10_brType(io_in_pds_10_brType),
    .io_in_pds_10_isRet(io_in_pds_10_isRet),
    .io_in_pds_11_isRVC(io_in_pds_11_isRVC),
    .io_in_pds_11_brType(io_in_pds_11_brType),
    .io_in_pds_11_isRet(io_in_pds_11_isRet),
    .io_in_pds_12_isRVC(io_in_pds_12_isRVC),
    .io_in_pds_12_brType(io_in_pds_12_brType),
    .io_in_pds_12_isRet(io_in_pds_12_isRet),
    .io_in_pds_13_isRVC(io_in_pds_13_isRVC),
    .io_in_pds_13_brType(io_in_pds_13_brType),
    .io_in_pds_13_isRet(io_in_pds_13_isRet),
    .io_in_pds_14_isRVC(io_in_pds_14_isRVC),
    .io_in_pds_14_brType(io_in_pds_14_brType),
    .io_in_pds_14_isRet(io_in_pds_14_isRet),
    .io_in_pds_15_isRVC(io_in_pds_15_isRVC),
    .io_in_pds_15_brType(io_in_pds_15_brType),
    .io_in_pds_15_isRet(io_in_pds_15_isRet),
    .io_in_pc_0(io_in_pc_0),
    .io_in_pc_1(io_in_pc_1),
    .io_in_pc_2(io_in_pc_2),
    .io_in_pc_3(io_in_pc_3),
    .io_in_pc_4(io_in_pc_4),
    .io_in_pc_5(io_in_pc_5),
    .io_in_pc_6(io_in_pc_6),
    .io_in_pc_7(io_in_pc_7),
    .io_in_pc_8(io_in_pc_8),
    .io_in_pc_9(io_in_pc_9),
    .io_in_pc_10(io_in_pc_10),
    .io_in_pc_11(io_in_pc_11),
    .io_in_pc_12(io_in_pc_12),
    .io_in_pc_13(io_in_pc_13),
    .io_in_pc_14(io_in_pc_14),
    .io_in_pc_15(io_in_pc_15),
    .io_in_fire_in(io_in_fire_in),
    .io_out_stage1Out_fixedRange_0(io_out_stage1Out_fixedRange_0),
    .io_out_stage1Out_fixedRange_1(io_out_stage1Out_fixedRange_1),
    .io_out_stage1Out_fixedRange_2(io_out_stage1Out_fixedRange_2),
    .io_out_stage1Out_fixedRange_3(io_out_stage1Out_fixedRange_3),
    .io_out_stage1Out_fixedRange_4(io_out_stage1Out_fixedRange_4),
    .io_out_stage1Out_fixedRange_5(io_out_stage1Out_fixedRange_5),
    .io_out_stage1Out_fixedRange_6(io_out_stage1Out_fixedRange_6),
    .io_out_stage1Out_fixedRange_7(io_out_stage1Out_fixedRange_7),
    .io_out_stage1Out_fixedRange_8(io_out_stage1Out_fixedRange_8),
    .io_out_stage1Out_fixedRange_9(io_out_stage1Out_fixedRange_9),
    .io_out_stage1Out_fixedRange_10(io_out_stage1Out_fixedRange_10),
    .io_out_stage1Out_fixedRange_11(io_out_stage1Out_fixedRange_11),
    .io_out_stage1Out_fixedRange_12(io_out_stage1Out_fixedRange_12),
    .io_out_stage1Out_fixedRange_13(io_out_stage1Out_fixedRange_13),
    .io_out_stage1Out_fixedRange_14(io_out_stage1Out_fixedRange_14),
    .io_out_stage1Out_fixedRange_15(io_out_stage1Out_fixedRange_15),
    .io_out_stage1Out_fixedTaken_0(io_out_stage1Out_fixedTaken_0),
    .io_out_stage1Out_fixedTaken_1(io_out_stage1Out_fixedTaken_1),
    .io_out_stage1Out_fixedTaken_2(io_out_stage1Out_fixedTaken_2),
    .io_out_stage1Out_fixedTaken_3(io_out_stage1Out_fixedTaken_3),
    .io_out_stage1Out_fixedTaken_4(io_out_stage1Out_fixedTaken_4),
    .io_out_stage1Out_fixedTaken_5(io_out_stage1Out_fixedTaken_5),
    .io_out_stage1Out_fixedTaken_6(io_out_stage1Out_fixedTaken_6),
    .io_out_stage1Out_fixedTaken_7(io_out_stage1Out_fixedTaken_7),
    .io_out_stage1Out_fixedTaken_8(io_out_stage1Out_fixedTaken_8),
    .io_out_stage1Out_fixedTaken_9(io_out_stage1Out_fixedTaken_9),
    .io_out_stage1Out_fixedTaken_10(io_out_stage1Out_fixedTaken_10),
    .io_out_stage1Out_fixedTaken_11(io_out_stage1Out_fixedTaken_11),
    .io_out_stage1Out_fixedTaken_12(io_out_stage1Out_fixedTaken_12),
    .io_out_stage1Out_fixedTaken_13(io_out_stage1Out_fixedTaken_13),
    .io_out_stage1Out_fixedTaken_14(io_out_stage1Out_fixedTaken_14),
    .io_out_stage1Out_fixedTaken_15(io_out_stage1Out_fixedTaken_15),
    .io_out_stage2Out_fixedTarget_0(io_out_stage2Out_fixedTarget_0),
    .io_out_stage2Out_fixedTarget_1(io_out_stage2Out_fixedTarget_1),
    .io_out_stage2Out_fixedTarget_2(io_out_stage2Out_fixedTarget_2),
    .io_out_stage2Out_fixedTarget_3(io_out_stage2Out_fixedTarget_3),
    .io_out_stage2Out_fixedTarget_4(io_out_stage2Out_fixedTarget_4),
    .io_out_stage2Out_fixedTarget_5(io_out_stage2Out_fixedTarget_5),
    .io_out_stage2Out_fixedTarget_6(io_out_stage2Out_fixedTarget_6),
    .io_out_stage2Out_fixedTarget_7(io_out_stage2Out_fixedTarget_7),
    .io_out_stage2Out_fixedTarget_8(io_out_stage2Out_fixedTarget_8),
    .io_out_stage2Out_fixedTarget_9(io_out_stage2Out_fixedTarget_9),
    .io_out_stage2Out_fixedTarget_10(io_out_stage2Out_fixedTarget_10),
    .io_out_stage2Out_fixedTarget_11(io_out_stage2Out_fixedTarget_11),
    .io_out_stage2Out_fixedTarget_12(io_out_stage2Out_fixedTarget_12),
    .io_out_stage2Out_fixedTarget_13(io_out_stage2Out_fixedTarget_13),
    .io_out_stage2Out_fixedTarget_14(io_out_stage2Out_fixedTarget_14),
    .io_out_stage2Out_fixedTarget_15(io_out_stage2Out_fixedTarget_15),
    .io_out_stage2Out_jalTarget_0(io_out_stage2Out_jalTarget_0),
    .io_out_stage2Out_jalTarget_1(io_out_stage2Out_jalTarget_1),
    .io_out_stage2Out_jalTarget_2(io_out_stage2Out_jalTarget_2),
    .io_out_stage2Out_jalTarget_3(io_out_stage2Out_jalTarget_3),
    .io_out_stage2Out_jalTarget_4(io_out_stage2Out_jalTarget_4),
    .io_out_stage2Out_jalTarget_5(io_out_stage2Out_jalTarget_5),
    .io_out_stage2Out_jalTarget_6(io_out_stage2Out_jalTarget_6),
    .io_out_stage2Out_jalTarget_7(io_out_stage2Out_jalTarget_7),
    .io_out_stage2Out_jalTarget_8(io_out_stage2Out_jalTarget_8),
    .io_out_stage2Out_jalTarget_9(io_out_stage2Out_jalTarget_9),
    .io_out_stage2Out_jalTarget_10(io_out_stage2Out_jalTarget_10),
    .io_out_stage2Out_jalTarget_11(io_out_stage2Out_jalTarget_11),
    .io_out_stage2Out_jalTarget_12(io_out_stage2Out_jalTarget_12),
    .io_out_stage2Out_jalTarget_13(io_out_stage2Out_jalTarget_13),
    .io_out_stage2Out_jalTarget_14(io_out_stage2Out_jalTarget_14),
    .io_out_stage2Out_jalTarget_15(io_out_stage2Out_jalTarget_15),
    .io_out_stage2Out_fixedMissPred_0(io_out_stage2Out_fixedMissPred_0),
    .io_out_stage2Out_fixedMissPred_1(io_out_stage2Out_fixedMissPred_1),
    .io_out_stage2Out_fixedMissPred_2(io_out_stage2Out_fixedMissPred_2),
    .io_out_stage2Out_fixedMissPred_3(io_out_stage2Out_fixedMissPred_3),
    .io_out_stage2Out_fixedMissPred_4(io_out_stage2Out_fixedMissPred_4),
    .io_out_stage2Out_fixedMissPred_5(io_out_stage2Out_fixedMissPred_5),
    .io_out_stage2Out_fixedMissPred_6(io_out_stage2Out_fixedMissPred_6),
    .io_out_stage2Out_fixedMissPred_7(io_out_stage2Out_fixedMissPred_7),
    .io_out_stage2Out_fixedMissPred_8(io_out_stage2Out_fixedMissPred_8),
    .io_out_stage2Out_fixedMissPred_9(io_out_stage2Out_fixedMissPred_9),
    .io_out_stage2Out_fixedMissPred_10(io_out_stage2Out_fixedMissPred_10),
    .io_out_stage2Out_fixedMissPred_11(io_out_stage2Out_fixedMissPred_11),
    .io_out_stage2Out_fixedMissPred_12(io_out_stage2Out_fixedMissPred_12),
    .io_out_stage2Out_fixedMissPred_13(io_out_stage2Out_fixedMissPred_13),
    .io_out_stage2Out_fixedMissPred_14(io_out_stage2Out_fixedMissPred_14),
    .io_out_stage2Out_fixedMissPred_15(io_out_stage2Out_fixedMissPred_15)
 );


endmodule

module F3Predecoder_top;

  wire [31:0] io_in_instr_0;
  wire [31:0] io_in_instr_1;
  wire [31:0] io_in_instr_2;
  wire [31:0] io_in_instr_3;
  wire [31:0] io_in_instr_4;
  wire [31:0] io_in_instr_5;
  wire [31:0] io_in_instr_6;
  wire [31:0] io_in_instr_7;
  wire [31:0] io_in_instr_8;
  wire [31:0] io_in_instr_9;
  wire [31:0] io_in_instr_10;
  wire [31:0] io_in_instr_11;
  wire [31:0] io_in_instr_12;
  wire [31:0] io_in_instr_13;
  wire [31:0] io_in_instr_14;
  wire [31:0] io_in_instr_15;
  wire [1:0] io_out_pd_0_brType;
  wire  io_out_pd_0_isCall;
  wire  io_out_pd_0_isRet;
  wire [1:0] io_out_pd_1_brType;
  wire  io_out_pd_1_isCall;
  wire  io_out_pd_1_isRet;
  wire [1:0] io_out_pd_2_brType;
  wire  io_out_pd_2_isCall;
  wire  io_out_pd_2_isRet;
  wire [1:0] io_out_pd_3_brType;
  wire  io_out_pd_3_isCall;
  wire  io_out_pd_3_isRet;
  wire [1:0] io_out_pd_4_brType;
  wire  io_out_pd_4_isCall;
  wire  io_out_pd_4_isRet;
  wire [1:0] io_out_pd_5_brType;
  wire  io_out_pd_5_isCall;
  wire  io_out_pd_5_isRet;
  wire [1:0] io_out_pd_6_brType;
  wire  io_out_pd_6_isCall;
  wire  io_out_pd_6_isRet;
  wire [1:0] io_out_pd_7_brType;
  wire  io_out_pd_7_isCall;
  wire  io_out_pd_7_isRet;
  wire [1:0] io_out_pd_8_brType;
  wire  io_out_pd_8_isCall;
  wire  io_out_pd_8_isRet;
  wire [1:0] io_out_pd_9_brType;
  wire  io_out_pd_9_isCall;
  wire  io_out_pd_9_isRet;
  wire [1:0] io_out_pd_10_brType;
  wire  io_out_pd_10_isCall;
  wire  io_out_pd_10_isRet;
  wire [1:0] io_out_pd_11_brType;
  wire  io_out_pd_11_isCall;
  wire  io_out_pd_11_isRet;
  wire [1:0] io_out_pd_12_brType;
  wire  io_out_pd_12_isCall;
  wire  io_out_pd_12_isRet;
  wire [1:0] io_out_pd_13_brType;
  wire  io_out_pd_13_isCall;
  wire  io_out_pd_13_isRet;
  wire [1:0] io_out_pd_14_brType;
  wire  io_out_pd_14_isCall;
  wire  io_out_pd_14_isRet;
  wire [1:0] io_out_pd_15_brType;
  wire  io_out_pd_15_isCall;
  wire  io_out_pd_15_isRet;


 F3Predecoder F3Predecoder(
    .io_in_instr_0(io_in_instr_0),
    .io_in_instr_1(io_in_instr_1),
    .io_in_instr_2(io_in_instr_2),
    .io_in_instr_3(io_in_instr_3),
    .io_in_instr_4(io_in_instr_4),
    .io_in_instr_5(io_in_instr_5),
    .io_in_instr_6(io_in_instr_6),
    .io_in_instr_7(io_in_instr_7),
    .io_in_instr_8(io_in_instr_8),
    .io_in_instr_9(io_in_instr_9),
    .io_in_instr_10(io_in_instr_10),
    .io_in_instr_11(io_in_instr_11),
    .io_in_instr_12(io_in_instr_12),
    .io_in_instr_13(io_in_instr_13),
    .io_in_instr_14(io_in_instr_14),
    .io_in_instr_15(io_in_instr_15),
    .io_out_pd_0_brType(io_out_pd_0_brType),
    .io_out_pd_0_isCall(io_out_pd_0_isCall),
    .io_out_pd_0_isRet(io_out_pd_0_isRet),
    .io_out_pd_1_brType(io_out_pd_1_brType),
    .io_out_pd_1_isCall(io_out_pd_1_isCall),
    .io_out_pd_1_isRet(io_out_pd_1_isRet),
    .io_out_pd_2_brType(io_out_pd_2_brType),
    .io_out_pd_2_isCall(io_out_pd_2_isCall),
    .io_out_pd_2_isRet(io_out_pd_2_isRet),
    .io_out_pd_3_brType(io_out_pd_3_brType),
    .io_out_pd_3_isCall(io_out_pd_3_isCall),
    .io_out_pd_3_isRet(io_out_pd_3_isRet),
    .io_out_pd_4_brType(io_out_pd_4_brType),
    .io_out_pd_4_isCall(io_out_pd_4_isCall),
    .io_out_pd_4_isRet(io_out_pd_4_isRet),
    .io_out_pd_5_brType(io_out_pd_5_brType),
    .io_out_pd_5_isCall(io_out_pd_5_isCall),
    .io_out_pd_5_isRet(io_out_pd_5_isRet),
    .io_out_pd_6_brType(io_out_pd_6_brType),
    .io_out_pd_6_isCall(io_out_pd_6_isCall),
    .io_out_pd_6_isRet(io_out_pd_6_isRet),
    .io_out_pd_7_brType(io_out_pd_7_brType),
    .io_out_pd_7_isCall(io_out_pd_7_isCall),
    .io_out_pd_7_isRet(io_out_pd_7_isRet),
    .io_out_pd_8_brType(io_out_pd_8_brType),
    .io_out_pd_8_isCall(io_out_pd_8_isCall),
    .io_out_pd_8_isRet(io_out_pd_8_isRet),
    .io_out_pd_9_brType(io_out_pd_9_brType),
    .io_out_pd_9_isCall(io_out_pd_9_isCall),
    .io_out_pd_9_isRet(io_out_pd_9_isRet),
    .io_out_pd_10_brType(io_out_pd_10_brType),
    .io_out_pd_10_isCall(io_out_pd_10_isCall),
    .io_out_pd_10_isRet(io_out_pd_10_isRet),
    .io_out_pd_11_brType(io_out_pd_11_brType),
    .io_out_pd_11_isCall(io_out_pd_11_isCall),
    .io_out_pd_11_isRet(io_out_pd_11_isRet),
    .io_out_pd_12_brType(io_out_pd_12_brType),
    .io_out_pd_12_isCall(io_out_pd_12_isCall),
    .io_out_pd_12_isRet(io_out_pd_12_isRet),
    .io_out_pd_13_brType(io_out_pd_13_brType),
    .io_out_pd_13_isCall(io_out_pd_13_isCall),
    .io_out_pd_13_isRet(io_out_pd_13_isRet),
    .io_out_pd_14_brType(io_out_pd_14_brType),
    .io_out_pd_14_isCall(io_out_pd_14_isCall),
    .io_out_pd_14_isRet(io_out_pd_14_isRet),
    .io_out_pd_15_brType(io_out_pd_15_brType),
    .io_out_pd_15_isCall(io_out_pd_15_isCall),
    .io_out_pd_15_isRet(io_out_pd_15_isRet)
 );


endmodule

module NewIFU_top;

  wire  clock;
  wire  reset;
  wire  io_ftqInter_fromFtq_req_ready;
  wire  io_ftqInter_fromFtq_req_valid;
  wire [49:0] io_ftqInter_fromFtq_req_bits_startAddr;
  wire [49:0] io_ftqInter_fromFtq_req_bits_nextlineStart;
  wire [49:0] io_ftqInter_fromFtq_req_bits_nextStartAddr;
  wire  io_ftqInter_fromFtq_req_bits_ftqIdx_flag;
  wire [5:0] io_ftqInter_fromFtq_req_bits_ftqIdx_value;
  wire  io_ftqInter_fromFtq_req_bits_ftqOffset_valid;
  wire [3:0] io_ftqInter_fromFtq_req_bits_ftqOffset_bits;
  wire  io_ftqInter_fromFtq_redirect_valid;
  wire  io_ftqInter_fromFtq_redirect_bits_ftqIdx_flag;
  wire [5:0] io_ftqInter_fromFtq_redirect_bits_ftqIdx_value;
  wire [3:0] io_ftqInter_fromFtq_redirect_bits_ftqOffset;
  wire  io_ftqInter_fromFtq_redirect_bits_level;
  wire  io_ftqInter_fromFtq_flushFromBpu_s2_valid;
  wire  io_ftqInter_fromFtq_flushFromBpu_s2_bits_flag;
  wire [5:0] io_ftqInter_fromFtq_flushFromBpu_s2_bits_value;
  wire  io_ftqInter_fromFtq_flushFromBpu_s3_valid;
  wire  io_ftqInter_fromFtq_flushFromBpu_s3_bits_flag;
  wire [5:0] io_ftqInter_fromFtq_flushFromBpu_s3_bits_value;
  wire  io_ftqInter_toFtq_pdWb_valid;
  wire [49:0] io_ftqInter_toFtq_pdWb_bits_pc_0;
  wire [49:0] io_ftqInter_toFtq_pdWb_bits_pc_1;
  wire [49:0] io_ftqInter_toFtq_pdWb_bits_pc_2;
  wire [49:0] io_ftqInter_toFtq_pdWb_bits_pc_3;
  wire [49:0] io_ftqInter_toFtq_pdWb_bits_pc_4;
  wire [49:0] io_ftqInter_toFtq_pdWb_bits_pc_5;
  wire [49:0] io_ftqInter_toFtq_pdWb_bits_pc_6;
  wire [49:0] io_ftqInter_toFtq_pdWb_bits_pc_7;
  wire [49:0] io_ftqInter_toFtq_pdWb_bits_pc_8;
  wire [49:0] io_ftqInter_toFtq_pdWb_bits_pc_9;
  wire [49:0] io_ftqInter_toFtq_pdWb_bits_pc_10;
  wire [49:0] io_ftqInter_toFtq_pdWb_bits_pc_11;
  wire [49:0] io_ftqInter_toFtq_pdWb_bits_pc_12;
  wire [49:0] io_ftqInter_toFtq_pdWb_bits_pc_13;
  wire [49:0] io_ftqInter_toFtq_pdWb_bits_pc_14;
  wire [49:0] io_ftqInter_toFtq_pdWb_bits_pc_15;
  wire  io_ftqInter_toFtq_pdWb_bits_pd_0_valid;
  wire  io_ftqInter_toFtq_pdWb_bits_pd_0_isRVC;
  wire [1:0] io_ftqInter_toFtq_pdWb_bits_pd_0_brType;
  wire  io_ftqInter_toFtq_pdWb_bits_pd_0_isCall;
  wire  io_ftqInter_toFtq_pdWb_bits_pd_0_isRet;
  wire  io_ftqInter_toFtq_pdWb_bits_pd_1_valid;
  wire  io_ftqInter_toFtq_pdWb_bits_pd_1_isRVC;
  wire [1:0] io_ftqInter_toFtq_pdWb_bits_pd_1_brType;
  wire  io_ftqInter_toFtq_pdWb_bits_pd_1_isCall;
  wire  io_ftqInter_toFtq_pdWb_bits_pd_1_isRet;
  wire  io_ftqInter_toFtq_pdWb_bits_pd_2_valid;
  wire  io_ftqInter_toFtq_pdWb_bits_pd_2_isRVC;
  wire [1:0] io_ftqInter_toFtq_pdWb_bits_pd_2_brType;
  wire  io_ftqInter_toFtq_pdWb_bits_pd_2_isCall;
  wire  io_ftqInter_toFtq_pdWb_bits_pd_2_isRet;
  wire  io_ftqInter_toFtq_pdWb_bits_pd_3_valid;
  wire  io_ftqInter_toFtq_pdWb_bits_pd_3_isRVC;
  wire [1:0] io_ftqInter_toFtq_pdWb_bits_pd_3_brType;
  wire  io_ftqInter_toFtq_pdWb_bits_pd_3_isCall;
  wire  io_ftqInter_toFtq_pdWb_bits_pd_3_isRet;
  wire  io_ftqInter_toFtq_pdWb_bits_pd_4_valid;
  wire  io_ftqInter_toFtq_pdWb_bits_pd_4_isRVC;
  wire [1:0] io_ftqInter_toFtq_pdWb_bits_pd_4_brType;
  wire  io_ftqInter_toFtq_pdWb_bits_pd_4_isCall;
  wire  io_ftqInter_toFtq_pdWb_bits_pd_4_isRet;
  wire  io_ftqInter_toFtq_pdWb_bits_pd_5_valid;
  wire  io_ftqInter_toFtq_pdWb_bits_pd_5_isRVC;
  wire [1:0] io_ftqInter_toFtq_pdWb_bits_pd_5_brType;
  wire  io_ftqInter_toFtq_pdWb_bits_pd_5_isCall;
  wire  io_ftqInter_toFtq_pdWb_bits_pd_5_isRet;
  wire  io_ftqInter_toFtq_pdWb_bits_pd_6_valid;
  wire  io_ftqInter_toFtq_pdWb_bits_pd_6_isRVC;
  wire [1:0] io_ftqInter_toFtq_pdWb_bits_pd_6_brType;
  wire  io_ftqInter_toFtq_pdWb_bits_pd_6_isCall;
  wire  io_ftqInter_toFtq_pdWb_bits_pd_6_isRet;
  wire  io_ftqInter_toFtq_pdWb_bits_pd_7_valid;
  wire  io_ftqInter_toFtq_pdWb_bits_pd_7_isRVC;
  wire [1:0] io_ftqInter_toFtq_pdWb_bits_pd_7_brType;
  wire  io_ftqInter_toFtq_pdWb_bits_pd_7_isCall;
  wire  io_ftqInter_toFtq_pdWb_bits_pd_7_isRet;
  wire  io_ftqInter_toFtq_pdWb_bits_pd_8_valid;
  wire  io_ftqInter_toFtq_pdWb_bits_pd_8_isRVC;
  wire [1:0] io_ftqInter_toFtq_pdWb_bits_pd_8_brType;
  wire  io_ftqInter_toFtq_pdWb_bits_pd_8_isCall;
  wire  io_ftqInter_toFtq_pdWb_bits_pd_8_isRet;
  wire  io_ftqInter_toFtq_pdWb_bits_pd_9_valid;
  wire  io_ftqInter_toFtq_pdWb_bits_pd_9_isRVC;
  wire [1:0] io_ftqInter_toFtq_pdWb_bits_pd_9_brType;
  wire  io_ftqInter_toFtq_pdWb_bits_pd_9_isCall;
  wire  io_ftqInter_toFtq_pdWb_bits_pd_9_isRet;
  wire  io_ftqInter_toFtq_pdWb_bits_pd_10_valid;
  wire  io_ftqInter_toFtq_pdWb_bits_pd_10_isRVC;
  wire [1:0] io_ftqInter_toFtq_pdWb_bits_pd_10_brType;
  wire  io_ftqInter_toFtq_pdWb_bits_pd_10_isCall;
  wire  io_ftqInter_toFtq_pdWb_bits_pd_10_isRet;
  wire  io_ftqInter_toFtq_pdWb_bits_pd_11_valid;
  wire  io_ftqInter_toFtq_pdWb_bits_pd_11_isRVC;
  wire [1:0] io_ftqInter_toFtq_pdWb_bits_pd_11_brType;
  wire  io_ftqInter_toFtq_pdWb_bits_pd_11_isCall;
  wire  io_ftqInter_toFtq_pdWb_bits_pd_11_isRet;
  wire  io_ftqInter_toFtq_pdWb_bits_pd_12_valid;
  wire  io_ftqInter_toFtq_pdWb_bits_pd_12_isRVC;
  wire [1:0] io_ftqInter_toFtq_pdWb_bits_pd_12_brType;
  wire  io_ftqInter_toFtq_pdWb_bits_pd_12_isCall;
  wire  io_ftqInter_toFtq_pdWb_bits_pd_12_isRet;
  wire  io_ftqInter_toFtq_pdWb_bits_pd_13_valid;
  wire  io_ftqInter_toFtq_pdWb_bits_pd_13_isRVC;
  wire [1:0] io_ftqInter_toFtq_pdWb_bits_pd_13_brType;
  wire  io_ftqInter_toFtq_pdWb_bits_pd_13_isCall;
  wire  io_ftqInter_toFtq_pdWb_bits_pd_13_isRet;
  wire  io_ftqInter_toFtq_pdWb_bits_pd_14_valid;
  wire  io_ftqInter_toFtq_pdWb_bits_pd_14_isRVC;
  wire [1:0] io_ftqInter_toFtq_pdWb_bits_pd_14_brType;
  wire  io_ftqInter_toFtq_pdWb_bits_pd_14_isCall;
  wire  io_ftqInter_toFtq_pdWb_bits_pd_14_isRet;
  wire  io_ftqInter_toFtq_pdWb_bits_pd_15_valid;
  wire  io_ftqInter_toFtq_pdWb_bits_pd_15_isRVC;
  wire [1:0] io_ftqInter_toFtq_pdWb_bits_pd_15_brType;
  wire  io_ftqInter_toFtq_pdWb_bits_pd_15_isCall;
  wire  io_ftqInter_toFtq_pdWb_bits_pd_15_isRet;
  wire  io_ftqInter_toFtq_pdWb_bits_ftqIdx_flag;
  wire [5:0] io_ftqInter_toFtq_pdWb_bits_ftqIdx_value;
  wire  io_ftqInter_toFtq_pdWb_bits_misOffset_valid;
  wire [3:0] io_ftqInter_toFtq_pdWb_bits_misOffset_bits;
  wire  io_ftqInter_toFtq_pdWb_bits_cfiOffset_valid;
  wire [49:0] io_ftqInter_toFtq_pdWb_bits_target;
  wire [49:0] io_ftqInter_toFtq_pdWb_bits_jalTarget;
  wire  io_ftqInter_toFtq_pdWb_bits_instrRange_0;
  wire  io_ftqInter_toFtq_pdWb_bits_instrRange_1;
  wire  io_ftqInter_toFtq_pdWb_bits_instrRange_2;
  wire  io_ftqInter_toFtq_pdWb_bits_instrRange_3;
  wire  io_ftqInter_toFtq_pdWb_bits_instrRange_4;
  wire  io_ftqInter_toFtq_pdWb_bits_instrRange_5;
  wire  io_ftqInter_toFtq_pdWb_bits_instrRange_6;
  wire  io_ftqInter_toFtq_pdWb_bits_instrRange_7;
  wire  io_ftqInter_toFtq_pdWb_bits_instrRange_8;
  wire  io_ftqInter_toFtq_pdWb_bits_instrRange_9;
  wire  io_ftqInter_toFtq_pdWb_bits_instrRange_10;
  wire  io_ftqInter_toFtq_pdWb_bits_instrRange_11;
  wire  io_ftqInter_toFtq_pdWb_bits_instrRange_12;
  wire  io_ftqInter_toFtq_pdWb_bits_instrRange_13;
  wire  io_ftqInter_toFtq_pdWb_bits_instrRange_14;
  wire  io_ftqInter_toFtq_pdWb_bits_instrRange_15;
  wire  io_icacheInter_icacheReady;
  wire  io_icacheInter_resp_valid;
  wire  io_icacheInter_resp_bits_doubleline;
  wire [49:0] io_icacheInter_resp_bits_vaddr_0;
  wire [49:0] io_icacheInter_resp_bits_vaddr_1;
  wire [511:0] io_icacheInter_resp_bits_data;
  wire [47:0] io_icacheInter_resp_bits_paddr_0;
  wire [1:0] io_icacheInter_resp_bits_exception_0;
  wire [1:0] io_icacheInter_resp_bits_exception_1;
  wire  io_icacheInter_resp_bits_pmp_mmio_0;
  wire  io_icacheInter_resp_bits_pmp_mmio_1;
  wire [1:0] io_icacheInter_resp_bits_itlb_pbmt_0;
  wire [1:0] io_icacheInter_resp_bits_itlb_pbmt_1;
  wire  io_icacheInter_resp_bits_backendException;
  wire [55:0] io_icacheInter_resp_bits_gpaddr;
  wire  io_icacheInter_resp_bits_isForVSnonLeafPTE;
  wire  io_icacheStop;
  wire  io_icachePerfInfo_only_0_hit;
  wire  io_icachePerfInfo_only_0_miss;
  wire  io_icachePerfInfo_hit_0_hit_1;
  wire  io_icachePerfInfo_hit_0_miss_1;
  wire  io_icachePerfInfo_miss_0_hit_1;
  wire  io_icachePerfInfo_miss_0_miss_1;
  wire  io_icachePerfInfo_bank_hit_1;
  wire  io_icachePerfInfo_hit;
  wire  io_toIbuffer_ready;
  wire  io_toIbuffer_valid;
  wire [31:0] io_toIbuffer_bits_instrs_0;
  wire [31:0] io_toIbuffer_bits_instrs_1;
  wire [31:0] io_toIbuffer_bits_instrs_2;
  wire [31:0] io_toIbuffer_bits_instrs_3;
  wire [31:0] io_toIbuffer_bits_instrs_4;
  wire [31:0] io_toIbuffer_bits_instrs_5;
  wire [31:0] io_toIbuffer_bits_instrs_6;
  wire [31:0] io_toIbuffer_bits_instrs_7;
  wire [31:0] io_toIbuffer_bits_instrs_8;
  wire [31:0] io_toIbuffer_bits_instrs_9;
  wire [31:0] io_toIbuffer_bits_instrs_10;
  wire [31:0] io_toIbuffer_bits_instrs_11;
  wire [31:0] io_toIbuffer_bits_instrs_12;
  wire [31:0] io_toIbuffer_bits_instrs_13;
  wire [31:0] io_toIbuffer_bits_instrs_14;
  wire [31:0] io_toIbuffer_bits_instrs_15;
  wire [15:0] io_toIbuffer_bits_valid;
  wire [15:0] io_toIbuffer_bits_enqEnable;
  wire  io_toIbuffer_bits_pd_0_isRVC;
  wire [1:0] io_toIbuffer_bits_pd_0_brType;
  wire  io_toIbuffer_bits_pd_1_isRVC;
  wire [1:0] io_toIbuffer_bits_pd_1_brType;
  wire  io_toIbuffer_bits_pd_2_isRVC;
  wire [1:0] io_toIbuffer_bits_pd_2_brType;
  wire  io_toIbuffer_bits_pd_3_isRVC;
  wire [1:0] io_toIbuffer_bits_pd_3_brType;
  wire  io_toIbuffer_bits_pd_4_isRVC;
  wire [1:0] io_toIbuffer_bits_pd_4_brType;
  wire  io_toIbuffer_bits_pd_5_isRVC;
  wire [1:0] io_toIbuffer_bits_pd_5_brType;
  wire  io_toIbuffer_bits_pd_6_isRVC;
  wire [1:0] io_toIbuffer_bits_pd_6_brType;
  wire  io_toIbuffer_bits_pd_7_isRVC;
  wire [1:0] io_toIbuffer_bits_pd_7_brType;
  wire  io_toIbuffer_bits_pd_8_isRVC;
  wire [1:0] io_toIbuffer_bits_pd_8_brType;
  wire  io_toIbuffer_bits_pd_9_isRVC;
  wire [1:0] io_toIbuffer_bits_pd_9_brType;
  wire  io_toIbuffer_bits_pd_10_isRVC;
  wire [1:0] io_toIbuffer_bits_pd_10_brType;
  wire  io_toIbuffer_bits_pd_11_isRVC;
  wire [1:0] io_toIbuffer_bits_pd_11_brType;
  wire  io_toIbuffer_bits_pd_12_isRVC;
  wire [1:0] io_toIbuffer_bits_pd_12_brType;
  wire  io_toIbuffer_bits_pd_13_isRVC;
  wire [1:0] io_toIbuffer_bits_pd_13_brType;
  wire  io_toIbuffer_bits_pd_14_isRVC;
  wire [1:0] io_toIbuffer_bits_pd_14_brType;
  wire  io_toIbuffer_bits_pd_15_isRVC;
  wire [1:0] io_toIbuffer_bits_pd_15_brType;
  wire [9:0] io_toIbuffer_bits_foldpc_0;
  wire [9:0] io_toIbuffer_bits_foldpc_1;
  wire [9:0] io_toIbuffer_bits_foldpc_2;
  wire [9:0] io_toIbuffer_bits_foldpc_3;
  wire [9:0] io_toIbuffer_bits_foldpc_4;
  wire [9:0] io_toIbuffer_bits_foldpc_5;
  wire [9:0] io_toIbuffer_bits_foldpc_6;
  wire [9:0] io_toIbuffer_bits_foldpc_7;
  wire [9:0] io_toIbuffer_bits_foldpc_8;
  wire [9:0] io_toIbuffer_bits_foldpc_9;
  wire [9:0] io_toIbuffer_bits_foldpc_10;
  wire [9:0] io_toIbuffer_bits_foldpc_11;
  wire [9:0] io_toIbuffer_bits_foldpc_12;
  wire [9:0] io_toIbuffer_bits_foldpc_13;
  wire [9:0] io_toIbuffer_bits_foldpc_14;
  wire [9:0] io_toIbuffer_bits_foldpc_15;
  wire  io_toIbuffer_bits_ftqOffset_0_valid;
  wire  io_toIbuffer_bits_ftqOffset_1_valid;
  wire  io_toIbuffer_bits_ftqOffset_2_valid;
  wire  io_toIbuffer_bits_ftqOffset_3_valid;
  wire  io_toIbuffer_bits_ftqOffset_4_valid;
  wire  io_toIbuffer_bits_ftqOffset_5_valid;
  wire  io_toIbuffer_bits_ftqOffset_6_valid;
  wire  io_toIbuffer_bits_ftqOffset_7_valid;
  wire  io_toIbuffer_bits_ftqOffset_8_valid;
  wire  io_toIbuffer_bits_ftqOffset_9_valid;
  wire  io_toIbuffer_bits_ftqOffset_10_valid;
  wire  io_toIbuffer_bits_ftqOffset_11_valid;
  wire  io_toIbuffer_bits_ftqOffset_12_valid;
  wire  io_toIbuffer_bits_ftqOffset_13_valid;
  wire  io_toIbuffer_bits_ftqOffset_14_valid;
  wire  io_toIbuffer_bits_ftqOffset_15_valid;
  wire  io_toIbuffer_bits_backendException_0;
  wire [1:0] io_toIbuffer_bits_exceptionType_0;
  wire [1:0] io_toIbuffer_bits_exceptionType_1;
  wire [1:0] io_toIbuffer_bits_exceptionType_2;
  wire [1:0] io_toIbuffer_bits_exceptionType_3;
  wire [1:0] io_toIbuffer_bits_exceptionType_4;
  wire [1:0] io_toIbuffer_bits_exceptionType_5;
  wire [1:0] io_toIbuffer_bits_exceptionType_6;
  wire [1:0] io_toIbuffer_bits_exceptionType_7;
  wire [1:0] io_toIbuffer_bits_exceptionType_8;
  wire [1:0] io_toIbuffer_bits_exceptionType_9;
  wire [1:0] io_toIbuffer_bits_exceptionType_10;
  wire [1:0] io_toIbuffer_bits_exceptionType_11;
  wire [1:0] io_toIbuffer_bits_exceptionType_12;
  wire [1:0] io_toIbuffer_bits_exceptionType_13;
  wire [1:0] io_toIbuffer_bits_exceptionType_14;
  wire [1:0] io_toIbuffer_bits_exceptionType_15;
  wire  io_toIbuffer_bits_crossPageIPFFix_0;
  wire  io_toIbuffer_bits_crossPageIPFFix_1;
  wire  io_toIbuffer_bits_crossPageIPFFix_2;
  wire  io_toIbuffer_bits_crossPageIPFFix_3;
  wire  io_toIbuffer_bits_crossPageIPFFix_4;
  wire  io_toIbuffer_bits_crossPageIPFFix_5;
  wire  io_toIbuffer_bits_crossPageIPFFix_6;
  wire  io_toIbuffer_bits_crossPageIPFFix_7;
  wire  io_toIbuffer_bits_crossPageIPFFix_8;
  wire  io_toIbuffer_bits_crossPageIPFFix_9;
  wire  io_toIbuffer_bits_crossPageIPFFix_10;
  wire  io_toIbuffer_bits_crossPageIPFFix_11;
  wire  io_toIbuffer_bits_crossPageIPFFix_12;
  wire  io_toIbuffer_bits_crossPageIPFFix_13;
  wire  io_toIbuffer_bits_crossPageIPFFix_14;
  wire  io_toIbuffer_bits_crossPageIPFFix_15;
  wire  io_toIbuffer_bits_illegalInstr_0;
  wire  io_toIbuffer_bits_illegalInstr_1;
  wire  io_toIbuffer_bits_illegalInstr_2;
  wire  io_toIbuffer_bits_illegalInstr_3;
  wire  io_toIbuffer_bits_illegalInstr_4;
  wire  io_toIbuffer_bits_illegalInstr_5;
  wire  io_toIbuffer_bits_illegalInstr_6;
  wire  io_toIbuffer_bits_illegalInstr_7;
  wire  io_toIbuffer_bits_illegalInstr_8;
  wire  io_toIbuffer_bits_illegalInstr_9;
  wire  io_toIbuffer_bits_illegalInstr_10;
  wire  io_toIbuffer_bits_illegalInstr_11;
  wire  io_toIbuffer_bits_illegalInstr_12;
  wire  io_toIbuffer_bits_illegalInstr_13;
  wire  io_toIbuffer_bits_illegalInstr_14;
  wire  io_toIbuffer_bits_illegalInstr_15;
  wire [3:0] io_toIbuffer_bits_triggered_0;
  wire [3:0] io_toIbuffer_bits_triggered_1;
  wire [3:0] io_toIbuffer_bits_triggered_2;
  wire [3:0] io_toIbuffer_bits_triggered_3;
  wire [3:0] io_toIbuffer_bits_triggered_4;
  wire [3:0] io_toIbuffer_bits_triggered_5;
  wire [3:0] io_toIbuffer_bits_triggered_6;
  wire [3:0] io_toIbuffer_bits_triggered_7;
  wire [3:0] io_toIbuffer_bits_triggered_8;
  wire [3:0] io_toIbuffer_bits_triggered_9;
  wire [3:0] io_toIbuffer_bits_triggered_10;
  wire [3:0] io_toIbuffer_bits_triggered_11;
  wire [3:0] io_toIbuffer_bits_triggered_12;
  wire [3:0] io_toIbuffer_bits_triggered_13;
  wire [3:0] io_toIbuffer_bits_triggered_14;
  wire [3:0] io_toIbuffer_bits_triggered_15;
  wire  io_toIbuffer_bits_isLastInFtqEntry_0;
  wire  io_toIbuffer_bits_isLastInFtqEntry_1;
  wire  io_toIbuffer_bits_isLastInFtqEntry_2;
  wire  io_toIbuffer_bits_isLastInFtqEntry_3;
  wire  io_toIbuffer_bits_isLastInFtqEntry_4;
  wire  io_toIbuffer_bits_isLastInFtqEntry_5;
  wire  io_toIbuffer_bits_isLastInFtqEntry_6;
  wire  io_toIbuffer_bits_isLastInFtqEntry_7;
  wire  io_toIbuffer_bits_isLastInFtqEntry_8;
  wire  io_toIbuffer_bits_isLastInFtqEntry_9;
  wire  io_toIbuffer_bits_isLastInFtqEntry_10;
  wire  io_toIbuffer_bits_isLastInFtqEntry_11;
  wire  io_toIbuffer_bits_isLastInFtqEntry_12;
  wire  io_toIbuffer_bits_isLastInFtqEntry_13;
  wire  io_toIbuffer_bits_isLastInFtqEntry_14;
  wire  io_toIbuffer_bits_isLastInFtqEntry_15;
  wire  io_toIbuffer_bits_ftqPtr_flag;
  wire [5:0] io_toIbuffer_bits_ftqPtr_value;
  wire  io_toBackend_gpaddrMem_wen;
  wire [5:0] io_toBackend_gpaddrMem_waddr;
  wire [55:0] io_toBackend_gpaddrMem_wdata_gpaddr;
  wire  io_toBackend_gpaddrMem_wdata_isForVSnonLeafPTE;
  wire  io_uncacheInter_fromUncache_valid;
  wire [31:0] io_uncacheInter_fromUncache_bits_data;
  wire  io_uncacheInter_toUncache_ready;
  wire  io_uncacheInter_toUncache_valid;
  wire [47:0] io_uncacheInter_toUncache_bits_addr;
  wire  io_frontendTrigger_tUpdate_valid;
  wire [1:0] io_frontendTrigger_tUpdate_bits_addr;
  wire [1:0] io_frontendTrigger_tUpdate_bits_tdata_matchType;
  wire  io_frontendTrigger_tUpdate_bits_tdata_select;
  wire [3:0] io_frontendTrigger_tUpdate_bits_tdata_action;
  wire  io_frontendTrigger_tUpdate_bits_tdata_chain;
  wire [63:0] io_frontendTrigger_tUpdate_bits_tdata_tdata2;
  wire  io_frontendTrigger_tEnableVec_0;
  wire  io_frontendTrigger_tEnableVec_1;
  wire  io_frontendTrigger_tEnableVec_2;
  wire  io_frontendTrigger_tEnableVec_3;
  wire  io_frontendTrigger_debugMode;
  wire  io_frontendTrigger_triggerCanRaiseBpExp;
  wire  io_rob_commits_0_valid;
  wire  io_rob_commits_0_bits_ftqIdx_flag;
  wire [5:0] io_rob_commits_0_bits_ftqIdx_value;
  wire [3:0] io_rob_commits_0_bits_ftqOffset;
  wire  io_rob_commits_1_valid;
  wire  io_rob_commits_1_bits_ftqIdx_flag;
  wire [5:0] io_rob_commits_1_bits_ftqIdx_value;
  wire [3:0] io_rob_commits_1_bits_ftqOffset;
  wire  io_rob_commits_2_valid;
  wire  io_rob_commits_2_bits_ftqIdx_flag;
  wire [5:0] io_rob_commits_2_bits_ftqIdx_value;
  wire [3:0] io_rob_commits_2_bits_ftqOffset;
  wire  io_rob_commits_3_valid;
  wire  io_rob_commits_3_bits_ftqIdx_flag;
  wire [5:0] io_rob_commits_3_bits_ftqIdx_value;
  wire [3:0] io_rob_commits_3_bits_ftqOffset;
  wire  io_rob_commits_4_valid;
  wire  io_rob_commits_4_bits_ftqIdx_flag;
  wire [5:0] io_rob_commits_4_bits_ftqIdx_value;
  wire [3:0] io_rob_commits_4_bits_ftqOffset;
  wire  io_rob_commits_5_valid;
  wire  io_rob_commits_5_bits_ftqIdx_flag;
  wire [5:0] io_rob_commits_5_bits_ftqIdx_value;
  wire [3:0] io_rob_commits_5_bits_ftqOffset;
  wire  io_rob_commits_6_valid;
  wire  io_rob_commits_6_bits_ftqIdx_flag;
  wire [5:0] io_rob_commits_6_bits_ftqIdx_value;
  wire [3:0] io_rob_commits_6_bits_ftqOffset;
  wire  io_rob_commits_7_valid;
  wire  io_rob_commits_7_bits_ftqIdx_flag;
  wire [5:0] io_rob_commits_7_bits_ftqIdx_value;
  wire [3:0] io_rob_commits_7_bits_ftqOffset;
  wire  io_iTLBInter_req_ready;
  wire  io_iTLBInter_req_valid;
  wire [49:0] io_iTLBInter_req_bits_vaddr;
  wire  io_iTLBInter_resp_ready;
  wire  io_iTLBInter_resp_valid;
  wire [47:0] io_iTLBInter_resp_bits_paddr_0;
  wire [63:0] io_iTLBInter_resp_bits_gpaddr_0;
  wire [1:0] io_iTLBInter_resp_bits_pbmt_0;
  wire  io_iTLBInter_resp_bits_isForVSnonLeafPTE;
  wire  io_iTLBInter_resp_bits_excp_0_gpf_instr;
  wire  io_iTLBInter_resp_bits_excp_0_pf_instr;
  wire  io_iTLBInter_resp_bits_excp_0_af_instr;
  wire [47:0] io_pmp_req_bits_addr;
  wire  io_pmp_resp_instr;
  wire  io_pmp_resp_mmio;
  wire  io_mmioCommitRead_mmioFtqPtr_flag;
  wire [5:0] io_mmioCommitRead_mmioFtqPtr_value;
  wire  io_mmioCommitRead_mmioLastCommit;
  wire  io_csr_fsIsOff;
  wire [5:0] io_perf_0_value;
  wire [5:0] io_perf_1_value;
  wire [5:0] io_perf_2_value;
  wire [5:0] io_perf_3_value;
  wire [5:0] io_perf_4_value;
  wire [5:0] io_perf_5_value;
  wire [5:0] io_perf_6_value;
  wire [5:0] io_perf_7_value;
  wire [5:0] io_perf_8_value;
  wire [5:0] io_perf_9_value;
  wire [5:0] io_perf_10_value;
  wire [5:0] io_perf_11_value;
  wire [5:0] io_perf_12_value;


 NewIFU NewIFU(
    .clock(clock),
    .reset(reset),
    .io_ftqInter_fromFtq_req_ready(io_ftqInter_fromFtq_req_ready),
    .io_ftqInter_fromFtq_req_valid(io_ftqInter_fromFtq_req_valid),
    .io_ftqInter_fromFtq_req_bits_startAddr(io_ftqInter_fromFtq_req_bits_startAddr),
    .io_ftqInter_fromFtq_req_bits_nextlineStart(io_ftqInter_fromFtq_req_bits_nextlineStart),
    .io_ftqInter_fromFtq_req_bits_nextStartAddr(io_ftqInter_fromFtq_req_bits_nextStartAddr),
    .io_ftqInter_fromFtq_req_bits_ftqIdx_flag(io_ftqInter_fromFtq_req_bits_ftqIdx_flag),
    .io_ftqInter_fromFtq_req_bits_ftqIdx_value(io_ftqInter_fromFtq_req_bits_ftqIdx_value),
    .io_ftqInter_fromFtq_req_bits_ftqOffset_valid(io_ftqInter_fromFtq_req_bits_ftqOffset_valid),
    .io_ftqInter_fromFtq_req_bits_ftqOffset_bits(io_ftqInter_fromFtq_req_bits_ftqOffset_bits),
    .io_ftqInter_fromFtq_redirect_valid(io_ftqInter_fromFtq_redirect_valid),
    .io_ftqInter_fromFtq_redirect_bits_ftqIdx_flag(io_ftqInter_fromFtq_redirect_bits_ftqIdx_flag),
    .io_ftqInter_fromFtq_redirect_bits_ftqIdx_value(io_ftqInter_fromFtq_redirect_bits_ftqIdx_value),
    .io_ftqInter_fromFtq_redirect_bits_ftqOffset(io_ftqInter_fromFtq_redirect_bits_ftqOffset),
    .io_ftqInter_fromFtq_redirect_bits_level(io_ftqInter_fromFtq_redirect_bits_level),
    .io_ftqInter_fromFtq_flushFromBpu_s2_valid(io_ftqInter_fromFtq_flushFromBpu_s2_valid),
    .io_ftqInter_fromFtq_flushFromBpu_s2_bits_flag(io_ftqInter_fromFtq_flushFromBpu_s2_bits_flag),
    .io_ftqInter_fromFtq_flushFromBpu_s2_bits_value(io_ftqInter_fromFtq_flushFromBpu_s2_bits_value),
    .io_ftqInter_fromFtq_flushFromBpu_s3_valid(io_ftqInter_fromFtq_flushFromBpu_s3_valid),
    .io_ftqInter_fromFtq_flushFromBpu_s3_bits_flag(io_ftqInter_fromFtq_flushFromBpu_s3_bits_flag),
    .io_ftqInter_fromFtq_flushFromBpu_s3_bits_value(io_ftqInter_fromFtq_flushFromBpu_s3_bits_value),
    .io_ftqInter_toFtq_pdWb_valid(io_ftqInter_toFtq_pdWb_valid),
    .io_ftqInter_toFtq_pdWb_bits_pc_0(io_ftqInter_toFtq_pdWb_bits_pc_0),
    .io_ftqInter_toFtq_pdWb_bits_pc_1(io_ftqInter_toFtq_pdWb_bits_pc_1),
    .io_ftqInter_toFtq_pdWb_bits_pc_2(io_ftqInter_toFtq_pdWb_bits_pc_2),
    .io_ftqInter_toFtq_pdWb_bits_pc_3(io_ftqInter_toFtq_pdWb_bits_pc_3),
    .io_ftqInter_toFtq_pdWb_bits_pc_4(io_ftqInter_toFtq_pdWb_bits_pc_4),
    .io_ftqInter_toFtq_pdWb_bits_pc_5(io_ftqInter_toFtq_pdWb_bits_pc_5),
    .io_ftqInter_toFtq_pdWb_bits_pc_6(io_ftqInter_toFtq_pdWb_bits_pc_6),
    .io_ftqInter_toFtq_pdWb_bits_pc_7(io_ftqInter_toFtq_pdWb_bits_pc_7),
    .io_ftqInter_toFtq_pdWb_bits_pc_8(io_ftqInter_toFtq_pdWb_bits_pc_8),
    .io_ftqInter_toFtq_pdWb_bits_pc_9(io_ftqInter_toFtq_pdWb_bits_pc_9),
    .io_ftqInter_toFtq_pdWb_bits_pc_10(io_ftqInter_toFtq_pdWb_bits_pc_10),
    .io_ftqInter_toFtq_pdWb_bits_pc_11(io_ftqInter_toFtq_pdWb_bits_pc_11),
    .io_ftqInter_toFtq_pdWb_bits_pc_12(io_ftqInter_toFtq_pdWb_bits_pc_12),
    .io_ftqInter_toFtq_pdWb_bits_pc_13(io_ftqInter_toFtq_pdWb_bits_pc_13),
    .io_ftqInter_toFtq_pdWb_bits_pc_14(io_ftqInter_toFtq_pdWb_bits_pc_14),
    .io_ftqInter_toFtq_pdWb_bits_pc_15(io_ftqInter_toFtq_pdWb_bits_pc_15),
    .io_ftqInter_toFtq_pdWb_bits_pd_0_valid(io_ftqInter_toFtq_pdWb_bits_pd_0_valid),
    .io_ftqInter_toFtq_pdWb_bits_pd_0_isRVC(io_ftqInter_toFtq_pdWb_bits_pd_0_isRVC),
    .io_ftqInter_toFtq_pdWb_bits_pd_0_brType(io_ftqInter_toFtq_pdWb_bits_pd_0_brType),
    .io_ftqInter_toFtq_pdWb_bits_pd_0_isCall(io_ftqInter_toFtq_pdWb_bits_pd_0_isCall),
    .io_ftqInter_toFtq_pdWb_bits_pd_0_isRet(io_ftqInter_toFtq_pdWb_bits_pd_0_isRet),
    .io_ftqInter_toFtq_pdWb_bits_pd_1_valid(io_ftqInter_toFtq_pdWb_bits_pd_1_valid),
    .io_ftqInter_toFtq_pdWb_bits_pd_1_isRVC(io_ftqInter_toFtq_pdWb_bits_pd_1_isRVC),
    .io_ftqInter_toFtq_pdWb_bits_pd_1_brType(io_ftqInter_toFtq_pdWb_bits_pd_1_brType),
    .io_ftqInter_toFtq_pdWb_bits_pd_1_isCall(io_ftqInter_toFtq_pdWb_bits_pd_1_isCall),
    .io_ftqInter_toFtq_pdWb_bits_pd_1_isRet(io_ftqInter_toFtq_pdWb_bits_pd_1_isRet),
    .io_ftqInter_toFtq_pdWb_bits_pd_2_valid(io_ftqInter_toFtq_pdWb_bits_pd_2_valid),
    .io_ftqInter_toFtq_pdWb_bits_pd_2_isRVC(io_ftqInter_toFtq_pdWb_bits_pd_2_isRVC),
    .io_ftqInter_toFtq_pdWb_bits_pd_2_brType(io_ftqInter_toFtq_pdWb_bits_pd_2_brType),
    .io_ftqInter_toFtq_pdWb_bits_pd_2_isCall(io_ftqInter_toFtq_pdWb_bits_pd_2_isCall),
    .io_ftqInter_toFtq_pdWb_bits_pd_2_isRet(io_ftqInter_toFtq_pdWb_bits_pd_2_isRet),
    .io_ftqInter_toFtq_pdWb_bits_pd_3_valid(io_ftqInter_toFtq_pdWb_bits_pd_3_valid),
    .io_ftqInter_toFtq_pdWb_bits_pd_3_isRVC(io_ftqInter_toFtq_pdWb_bits_pd_3_isRVC),
    .io_ftqInter_toFtq_pdWb_bits_pd_3_brType(io_ftqInter_toFtq_pdWb_bits_pd_3_brType),
    .io_ftqInter_toFtq_pdWb_bits_pd_3_isCall(io_ftqInter_toFtq_pdWb_bits_pd_3_isCall),
    .io_ftqInter_toFtq_pdWb_bits_pd_3_isRet(io_ftqInter_toFtq_pdWb_bits_pd_3_isRet),
    .io_ftqInter_toFtq_pdWb_bits_pd_4_valid(io_ftqInter_toFtq_pdWb_bits_pd_4_valid),
    .io_ftqInter_toFtq_pdWb_bits_pd_4_isRVC(io_ftqInter_toFtq_pdWb_bits_pd_4_isRVC),
    .io_ftqInter_toFtq_pdWb_bits_pd_4_brType(io_ftqInter_toFtq_pdWb_bits_pd_4_brType),
    .io_ftqInter_toFtq_pdWb_bits_pd_4_isCall(io_ftqInter_toFtq_pdWb_bits_pd_4_isCall),
    .io_ftqInter_toFtq_pdWb_bits_pd_4_isRet(io_ftqInter_toFtq_pdWb_bits_pd_4_isRet),
    .io_ftqInter_toFtq_pdWb_bits_pd_5_valid(io_ftqInter_toFtq_pdWb_bits_pd_5_valid),
    .io_ftqInter_toFtq_pdWb_bits_pd_5_isRVC(io_ftqInter_toFtq_pdWb_bits_pd_5_isRVC),
    .io_ftqInter_toFtq_pdWb_bits_pd_5_brType(io_ftqInter_toFtq_pdWb_bits_pd_5_brType),
    .io_ftqInter_toFtq_pdWb_bits_pd_5_isCall(io_ftqInter_toFtq_pdWb_bits_pd_5_isCall),
    .io_ftqInter_toFtq_pdWb_bits_pd_5_isRet(io_ftqInter_toFtq_pdWb_bits_pd_5_isRet),
    .io_ftqInter_toFtq_pdWb_bits_pd_6_valid(io_ftqInter_toFtq_pdWb_bits_pd_6_valid),
    .io_ftqInter_toFtq_pdWb_bits_pd_6_isRVC(io_ftqInter_toFtq_pdWb_bits_pd_6_isRVC),
    .io_ftqInter_toFtq_pdWb_bits_pd_6_brType(io_ftqInter_toFtq_pdWb_bits_pd_6_brType),
    .io_ftqInter_toFtq_pdWb_bits_pd_6_isCall(io_ftqInter_toFtq_pdWb_bits_pd_6_isCall),
    .io_ftqInter_toFtq_pdWb_bits_pd_6_isRet(io_ftqInter_toFtq_pdWb_bits_pd_6_isRet),
    .io_ftqInter_toFtq_pdWb_bits_pd_7_valid(io_ftqInter_toFtq_pdWb_bits_pd_7_valid),
    .io_ftqInter_toFtq_pdWb_bits_pd_7_isRVC(io_ftqInter_toFtq_pdWb_bits_pd_7_isRVC),
    .io_ftqInter_toFtq_pdWb_bits_pd_7_brType(io_ftqInter_toFtq_pdWb_bits_pd_7_brType),
    .io_ftqInter_toFtq_pdWb_bits_pd_7_isCall(io_ftqInter_toFtq_pdWb_bits_pd_7_isCall),
    .io_ftqInter_toFtq_pdWb_bits_pd_7_isRet(io_ftqInter_toFtq_pdWb_bits_pd_7_isRet),
    .io_ftqInter_toFtq_pdWb_bits_pd_8_valid(io_ftqInter_toFtq_pdWb_bits_pd_8_valid),
    .io_ftqInter_toFtq_pdWb_bits_pd_8_isRVC(io_ftqInter_toFtq_pdWb_bits_pd_8_isRVC),
    .io_ftqInter_toFtq_pdWb_bits_pd_8_brType(io_ftqInter_toFtq_pdWb_bits_pd_8_brType),
    .io_ftqInter_toFtq_pdWb_bits_pd_8_isCall(io_ftqInter_toFtq_pdWb_bits_pd_8_isCall),
    .io_ftqInter_toFtq_pdWb_bits_pd_8_isRet(io_ftqInter_toFtq_pdWb_bits_pd_8_isRet),
    .io_ftqInter_toFtq_pdWb_bits_pd_9_valid(io_ftqInter_toFtq_pdWb_bits_pd_9_valid),
    .io_ftqInter_toFtq_pdWb_bits_pd_9_isRVC(io_ftqInter_toFtq_pdWb_bits_pd_9_isRVC),
    .io_ftqInter_toFtq_pdWb_bits_pd_9_brType(io_ftqInter_toFtq_pdWb_bits_pd_9_brType),
    .io_ftqInter_toFtq_pdWb_bits_pd_9_isCall(io_ftqInter_toFtq_pdWb_bits_pd_9_isCall),
    .io_ftqInter_toFtq_pdWb_bits_pd_9_isRet(io_ftqInter_toFtq_pdWb_bits_pd_9_isRet),
    .io_ftqInter_toFtq_pdWb_bits_pd_10_valid(io_ftqInter_toFtq_pdWb_bits_pd_10_valid),
    .io_ftqInter_toFtq_pdWb_bits_pd_10_isRVC(io_ftqInter_toFtq_pdWb_bits_pd_10_isRVC),
    .io_ftqInter_toFtq_pdWb_bits_pd_10_brType(io_ftqInter_toFtq_pdWb_bits_pd_10_brType),
    .io_ftqInter_toFtq_pdWb_bits_pd_10_isCall(io_ftqInter_toFtq_pdWb_bits_pd_10_isCall),
    .io_ftqInter_toFtq_pdWb_bits_pd_10_isRet(io_ftqInter_toFtq_pdWb_bits_pd_10_isRet),
    .io_ftqInter_toFtq_pdWb_bits_pd_11_valid(io_ftqInter_toFtq_pdWb_bits_pd_11_valid),
    .io_ftqInter_toFtq_pdWb_bits_pd_11_isRVC(io_ftqInter_toFtq_pdWb_bits_pd_11_isRVC),
    .io_ftqInter_toFtq_pdWb_bits_pd_11_brType(io_ftqInter_toFtq_pdWb_bits_pd_11_brType),
    .io_ftqInter_toFtq_pdWb_bits_pd_11_isCall(io_ftqInter_toFtq_pdWb_bits_pd_11_isCall),
    .io_ftqInter_toFtq_pdWb_bits_pd_11_isRet(io_ftqInter_toFtq_pdWb_bits_pd_11_isRet),
    .io_ftqInter_toFtq_pdWb_bits_pd_12_valid(io_ftqInter_toFtq_pdWb_bits_pd_12_valid),
    .io_ftqInter_toFtq_pdWb_bits_pd_12_isRVC(io_ftqInter_toFtq_pdWb_bits_pd_12_isRVC),
    .io_ftqInter_toFtq_pdWb_bits_pd_12_brType(io_ftqInter_toFtq_pdWb_bits_pd_12_brType),
    .io_ftqInter_toFtq_pdWb_bits_pd_12_isCall(io_ftqInter_toFtq_pdWb_bits_pd_12_isCall),
    .io_ftqInter_toFtq_pdWb_bits_pd_12_isRet(io_ftqInter_toFtq_pdWb_bits_pd_12_isRet),
    .io_ftqInter_toFtq_pdWb_bits_pd_13_valid(io_ftqInter_toFtq_pdWb_bits_pd_13_valid),
    .io_ftqInter_toFtq_pdWb_bits_pd_13_isRVC(io_ftqInter_toFtq_pdWb_bits_pd_13_isRVC),
    .io_ftqInter_toFtq_pdWb_bits_pd_13_brType(io_ftqInter_toFtq_pdWb_bits_pd_13_brType),
    .io_ftqInter_toFtq_pdWb_bits_pd_13_isCall(io_ftqInter_toFtq_pdWb_bits_pd_13_isCall),
    .io_ftqInter_toFtq_pdWb_bits_pd_13_isRet(io_ftqInter_toFtq_pdWb_bits_pd_13_isRet),
    .io_ftqInter_toFtq_pdWb_bits_pd_14_valid(io_ftqInter_toFtq_pdWb_bits_pd_14_valid),
    .io_ftqInter_toFtq_pdWb_bits_pd_14_isRVC(io_ftqInter_toFtq_pdWb_bits_pd_14_isRVC),
    .io_ftqInter_toFtq_pdWb_bits_pd_14_brType(io_ftqInter_toFtq_pdWb_bits_pd_14_brType),
    .io_ftqInter_toFtq_pdWb_bits_pd_14_isCall(io_ftqInter_toFtq_pdWb_bits_pd_14_isCall),
    .io_ftqInter_toFtq_pdWb_bits_pd_14_isRet(io_ftqInter_toFtq_pdWb_bits_pd_14_isRet),
    .io_ftqInter_toFtq_pdWb_bits_pd_15_valid(io_ftqInter_toFtq_pdWb_bits_pd_15_valid),
    .io_ftqInter_toFtq_pdWb_bits_pd_15_isRVC(io_ftqInter_toFtq_pdWb_bits_pd_15_isRVC),
    .io_ftqInter_toFtq_pdWb_bits_pd_15_brType(io_ftqInter_toFtq_pdWb_bits_pd_15_brType),
    .io_ftqInter_toFtq_pdWb_bits_pd_15_isCall(io_ftqInter_toFtq_pdWb_bits_pd_15_isCall),
    .io_ftqInter_toFtq_pdWb_bits_pd_15_isRet(io_ftqInter_toFtq_pdWb_bits_pd_15_isRet),
    .io_ftqInter_toFtq_pdWb_bits_ftqIdx_flag(io_ftqInter_toFtq_pdWb_bits_ftqIdx_flag),
    .io_ftqInter_toFtq_pdWb_bits_ftqIdx_value(io_ftqInter_toFtq_pdWb_bits_ftqIdx_value),
    .io_ftqInter_toFtq_pdWb_bits_misOffset_valid(io_ftqInter_toFtq_pdWb_bits_misOffset_valid),
    .io_ftqInter_toFtq_pdWb_bits_misOffset_bits(io_ftqInter_toFtq_pdWb_bits_misOffset_bits),
    .io_ftqInter_toFtq_pdWb_bits_cfiOffset_valid(io_ftqInter_toFtq_pdWb_bits_cfiOffset_valid),
    .io_ftqInter_toFtq_pdWb_bits_target(io_ftqInter_toFtq_pdWb_bits_target),
    .io_ftqInter_toFtq_pdWb_bits_jalTarget(io_ftqInter_toFtq_pdWb_bits_jalTarget),
    .io_ftqInter_toFtq_pdWb_bits_instrRange_0(io_ftqInter_toFtq_pdWb_bits_instrRange_0),
    .io_ftqInter_toFtq_pdWb_bits_instrRange_1(io_ftqInter_toFtq_pdWb_bits_instrRange_1),
    .io_ftqInter_toFtq_pdWb_bits_instrRange_2(io_ftqInter_toFtq_pdWb_bits_instrRange_2),
    .io_ftqInter_toFtq_pdWb_bits_instrRange_3(io_ftqInter_toFtq_pdWb_bits_instrRange_3),
    .io_ftqInter_toFtq_pdWb_bits_instrRange_4(io_ftqInter_toFtq_pdWb_bits_instrRange_4),
    .io_ftqInter_toFtq_pdWb_bits_instrRange_5(io_ftqInter_toFtq_pdWb_bits_instrRange_5),
    .io_ftqInter_toFtq_pdWb_bits_instrRange_6(io_ftqInter_toFtq_pdWb_bits_instrRange_6),
    .io_ftqInter_toFtq_pdWb_bits_instrRange_7(io_ftqInter_toFtq_pdWb_bits_instrRange_7),
    .io_ftqInter_toFtq_pdWb_bits_instrRange_8(io_ftqInter_toFtq_pdWb_bits_instrRange_8),
    .io_ftqInter_toFtq_pdWb_bits_instrRange_9(io_ftqInter_toFtq_pdWb_bits_instrRange_9),
    .io_ftqInter_toFtq_pdWb_bits_instrRange_10(io_ftqInter_toFtq_pdWb_bits_instrRange_10),
    .io_ftqInter_toFtq_pdWb_bits_instrRange_11(io_ftqInter_toFtq_pdWb_bits_instrRange_11),
    .io_ftqInter_toFtq_pdWb_bits_instrRange_12(io_ftqInter_toFtq_pdWb_bits_instrRange_12),
    .io_ftqInter_toFtq_pdWb_bits_instrRange_13(io_ftqInter_toFtq_pdWb_bits_instrRange_13),
    .io_ftqInter_toFtq_pdWb_bits_instrRange_14(io_ftqInter_toFtq_pdWb_bits_instrRange_14),
    .io_ftqInter_toFtq_pdWb_bits_instrRange_15(io_ftqInter_toFtq_pdWb_bits_instrRange_15),
    .io_icacheInter_icacheReady(io_icacheInter_icacheReady),
    .io_icacheInter_resp_valid(io_icacheInter_resp_valid),
    .io_icacheInter_resp_bits_doubleline(io_icacheInter_resp_bits_doubleline),
    .io_icacheInter_resp_bits_vaddr_0(io_icacheInter_resp_bits_vaddr_0),
    .io_icacheInter_resp_bits_vaddr_1(io_icacheInter_resp_bits_vaddr_1),
    .io_icacheInter_resp_bits_data(io_icacheInter_resp_bits_data),
    .io_icacheInter_resp_bits_paddr_0(io_icacheInter_resp_bits_paddr_0),
    .io_icacheInter_resp_bits_exception_0(io_icacheInter_resp_bits_exception_0),
    .io_icacheInter_resp_bits_exception_1(io_icacheInter_resp_bits_exception_1),
    .io_icacheInter_resp_bits_pmp_mmio_0(io_icacheInter_resp_bits_pmp_mmio_0),
    .io_icacheInter_resp_bits_pmp_mmio_1(io_icacheInter_resp_bits_pmp_mmio_1),
    .io_icacheInter_resp_bits_itlb_pbmt_0(io_icacheInter_resp_bits_itlb_pbmt_0),
    .io_icacheInter_resp_bits_itlb_pbmt_1(io_icacheInter_resp_bits_itlb_pbmt_1),
    .io_icacheInter_resp_bits_backendException(io_icacheInter_resp_bits_backendException),
    .io_icacheInter_resp_bits_gpaddr(io_icacheInter_resp_bits_gpaddr),
    .io_icacheInter_resp_bits_isForVSnonLeafPTE(io_icacheInter_resp_bits_isForVSnonLeafPTE),
    .io_icacheStop(io_icacheStop),
    .io_icachePerfInfo_only_0_hit(io_icachePerfInfo_only_0_hit),
    .io_icachePerfInfo_only_0_miss(io_icachePerfInfo_only_0_miss),
    .io_icachePerfInfo_hit_0_hit_1(io_icachePerfInfo_hit_0_hit_1),
    .io_icachePerfInfo_hit_0_miss_1(io_icachePerfInfo_hit_0_miss_1),
    .io_icachePerfInfo_miss_0_hit_1(io_icachePerfInfo_miss_0_hit_1),
    .io_icachePerfInfo_miss_0_miss_1(io_icachePerfInfo_miss_0_miss_1),
    .io_icachePerfInfo_bank_hit_1(io_icachePerfInfo_bank_hit_1),
    .io_icachePerfInfo_hit(io_icachePerfInfo_hit),
    .io_toIbuffer_ready(io_toIbuffer_ready),
    .io_toIbuffer_valid(io_toIbuffer_valid),
    .io_toIbuffer_bits_instrs_0(io_toIbuffer_bits_instrs_0),
    .io_toIbuffer_bits_instrs_1(io_toIbuffer_bits_instrs_1),
    .io_toIbuffer_bits_instrs_2(io_toIbuffer_bits_instrs_2),
    .io_toIbuffer_bits_instrs_3(io_toIbuffer_bits_instrs_3),
    .io_toIbuffer_bits_instrs_4(io_toIbuffer_bits_instrs_4),
    .io_toIbuffer_bits_instrs_5(io_toIbuffer_bits_instrs_5),
    .io_toIbuffer_bits_instrs_6(io_toIbuffer_bits_instrs_6),
    .io_toIbuffer_bits_instrs_7(io_toIbuffer_bits_instrs_7),
    .io_toIbuffer_bits_instrs_8(io_toIbuffer_bits_instrs_8),
    .io_toIbuffer_bits_instrs_9(io_toIbuffer_bits_instrs_9),
    .io_toIbuffer_bits_instrs_10(io_toIbuffer_bits_instrs_10),
    .io_toIbuffer_bits_instrs_11(io_toIbuffer_bits_instrs_11),
    .io_toIbuffer_bits_instrs_12(io_toIbuffer_bits_instrs_12),
    .io_toIbuffer_bits_instrs_13(io_toIbuffer_bits_instrs_13),
    .io_toIbuffer_bits_instrs_14(io_toIbuffer_bits_instrs_14),
    .io_toIbuffer_bits_instrs_15(io_toIbuffer_bits_instrs_15),
    .io_toIbuffer_bits_valid(io_toIbuffer_bits_valid),
    .io_toIbuffer_bits_enqEnable(io_toIbuffer_bits_enqEnable),
    .io_toIbuffer_bits_pd_0_isRVC(io_toIbuffer_bits_pd_0_isRVC),
    .io_toIbuffer_bits_pd_0_brType(io_toIbuffer_bits_pd_0_brType),
    .io_toIbuffer_bits_pd_1_isRVC(io_toIbuffer_bits_pd_1_isRVC),
    .io_toIbuffer_bits_pd_1_brType(io_toIbuffer_bits_pd_1_brType),
    .io_toIbuffer_bits_pd_2_isRVC(io_toIbuffer_bits_pd_2_isRVC),
    .io_toIbuffer_bits_pd_2_brType(io_toIbuffer_bits_pd_2_brType),
    .io_toIbuffer_bits_pd_3_isRVC(io_toIbuffer_bits_pd_3_isRVC),
    .io_toIbuffer_bits_pd_3_brType(io_toIbuffer_bits_pd_3_brType),
    .io_toIbuffer_bits_pd_4_isRVC(io_toIbuffer_bits_pd_4_isRVC),
    .io_toIbuffer_bits_pd_4_brType(io_toIbuffer_bits_pd_4_brType),
    .io_toIbuffer_bits_pd_5_isRVC(io_toIbuffer_bits_pd_5_isRVC),
    .io_toIbuffer_bits_pd_5_brType(io_toIbuffer_bits_pd_5_brType),
    .io_toIbuffer_bits_pd_6_isRVC(io_toIbuffer_bits_pd_6_isRVC),
    .io_toIbuffer_bits_pd_6_brType(io_toIbuffer_bits_pd_6_brType),
    .io_toIbuffer_bits_pd_7_isRVC(io_toIbuffer_bits_pd_7_isRVC),
    .io_toIbuffer_bits_pd_7_brType(io_toIbuffer_bits_pd_7_brType),
    .io_toIbuffer_bits_pd_8_isRVC(io_toIbuffer_bits_pd_8_isRVC),
    .io_toIbuffer_bits_pd_8_brType(io_toIbuffer_bits_pd_8_brType),
    .io_toIbuffer_bits_pd_9_isRVC(io_toIbuffer_bits_pd_9_isRVC),
    .io_toIbuffer_bits_pd_9_brType(io_toIbuffer_bits_pd_9_brType),
    .io_toIbuffer_bits_pd_10_isRVC(io_toIbuffer_bits_pd_10_isRVC),
    .io_toIbuffer_bits_pd_10_brType(io_toIbuffer_bits_pd_10_brType),
    .io_toIbuffer_bits_pd_11_isRVC(io_toIbuffer_bits_pd_11_isRVC),
    .io_toIbuffer_bits_pd_11_brType(io_toIbuffer_bits_pd_11_brType),
    .io_toIbuffer_bits_pd_12_isRVC(io_toIbuffer_bits_pd_12_isRVC),
    .io_toIbuffer_bits_pd_12_brType(io_toIbuffer_bits_pd_12_brType),
    .io_toIbuffer_bits_pd_13_isRVC(io_toIbuffer_bits_pd_13_isRVC),
    .io_toIbuffer_bits_pd_13_brType(io_toIbuffer_bits_pd_13_brType),
    .io_toIbuffer_bits_pd_14_isRVC(io_toIbuffer_bits_pd_14_isRVC),
    .io_toIbuffer_bits_pd_14_brType(io_toIbuffer_bits_pd_14_brType),
    .io_toIbuffer_bits_pd_15_isRVC(io_toIbuffer_bits_pd_15_isRVC),
    .io_toIbuffer_bits_pd_15_brType(io_toIbuffer_bits_pd_15_brType),
    .io_toIbuffer_bits_foldpc_0(io_toIbuffer_bits_foldpc_0),
    .io_toIbuffer_bits_foldpc_1(io_toIbuffer_bits_foldpc_1),
    .io_toIbuffer_bits_foldpc_2(io_toIbuffer_bits_foldpc_2),
    .io_toIbuffer_bits_foldpc_3(io_toIbuffer_bits_foldpc_3),
    .io_toIbuffer_bits_foldpc_4(io_toIbuffer_bits_foldpc_4),
    .io_toIbuffer_bits_foldpc_5(io_toIbuffer_bits_foldpc_5),
    .io_toIbuffer_bits_foldpc_6(io_toIbuffer_bits_foldpc_6),
    .io_toIbuffer_bits_foldpc_7(io_toIbuffer_bits_foldpc_7),
    .io_toIbuffer_bits_foldpc_8(io_toIbuffer_bits_foldpc_8),
    .io_toIbuffer_bits_foldpc_9(io_toIbuffer_bits_foldpc_9),
    .io_toIbuffer_bits_foldpc_10(io_toIbuffer_bits_foldpc_10),
    .io_toIbuffer_bits_foldpc_11(io_toIbuffer_bits_foldpc_11),
    .io_toIbuffer_bits_foldpc_12(io_toIbuffer_bits_foldpc_12),
    .io_toIbuffer_bits_foldpc_13(io_toIbuffer_bits_foldpc_13),
    .io_toIbuffer_bits_foldpc_14(io_toIbuffer_bits_foldpc_14),
    .io_toIbuffer_bits_foldpc_15(io_toIbuffer_bits_foldpc_15),
    .io_toIbuffer_bits_ftqOffset_0_valid(io_toIbuffer_bits_ftqOffset_0_valid),
    .io_toIbuffer_bits_ftqOffset_1_valid(io_toIbuffer_bits_ftqOffset_1_valid),
    .io_toIbuffer_bits_ftqOffset_2_valid(io_toIbuffer_bits_ftqOffset_2_valid),
    .io_toIbuffer_bits_ftqOffset_3_valid(io_toIbuffer_bits_ftqOffset_3_valid),
    .io_toIbuffer_bits_ftqOffset_4_valid(io_toIbuffer_bits_ftqOffset_4_valid),
    .io_toIbuffer_bits_ftqOffset_5_valid(io_toIbuffer_bits_ftqOffset_5_valid),
    .io_toIbuffer_bits_ftqOffset_6_valid(io_toIbuffer_bits_ftqOffset_6_valid),
    .io_toIbuffer_bits_ftqOffset_7_valid(io_toIbuffer_bits_ftqOffset_7_valid),
    .io_toIbuffer_bits_ftqOffset_8_valid(io_toIbuffer_bits_ftqOffset_8_valid),
    .io_toIbuffer_bits_ftqOffset_9_valid(io_toIbuffer_bits_ftqOffset_9_valid),
    .io_toIbuffer_bits_ftqOffset_10_valid(io_toIbuffer_bits_ftqOffset_10_valid),
    .io_toIbuffer_bits_ftqOffset_11_valid(io_toIbuffer_bits_ftqOffset_11_valid),
    .io_toIbuffer_bits_ftqOffset_12_valid(io_toIbuffer_bits_ftqOffset_12_valid),
    .io_toIbuffer_bits_ftqOffset_13_valid(io_toIbuffer_bits_ftqOffset_13_valid),
    .io_toIbuffer_bits_ftqOffset_14_valid(io_toIbuffer_bits_ftqOffset_14_valid),
    .io_toIbuffer_bits_ftqOffset_15_valid(io_toIbuffer_bits_ftqOffset_15_valid),
    .io_toIbuffer_bits_backendException_0(io_toIbuffer_bits_backendException_0),
    .io_toIbuffer_bits_exceptionType_0(io_toIbuffer_bits_exceptionType_0),
    .io_toIbuffer_bits_exceptionType_1(io_toIbuffer_bits_exceptionType_1),
    .io_toIbuffer_bits_exceptionType_2(io_toIbuffer_bits_exceptionType_2),
    .io_toIbuffer_bits_exceptionType_3(io_toIbuffer_bits_exceptionType_3),
    .io_toIbuffer_bits_exceptionType_4(io_toIbuffer_bits_exceptionType_4),
    .io_toIbuffer_bits_exceptionType_5(io_toIbuffer_bits_exceptionType_5),
    .io_toIbuffer_bits_exceptionType_6(io_toIbuffer_bits_exceptionType_6),
    .io_toIbuffer_bits_exceptionType_7(io_toIbuffer_bits_exceptionType_7),
    .io_toIbuffer_bits_exceptionType_8(io_toIbuffer_bits_exceptionType_8),
    .io_toIbuffer_bits_exceptionType_9(io_toIbuffer_bits_exceptionType_9),
    .io_toIbuffer_bits_exceptionType_10(io_toIbuffer_bits_exceptionType_10),
    .io_toIbuffer_bits_exceptionType_11(io_toIbuffer_bits_exceptionType_11),
    .io_toIbuffer_bits_exceptionType_12(io_toIbuffer_bits_exceptionType_12),
    .io_toIbuffer_bits_exceptionType_13(io_toIbuffer_bits_exceptionType_13),
    .io_toIbuffer_bits_exceptionType_14(io_toIbuffer_bits_exceptionType_14),
    .io_toIbuffer_bits_exceptionType_15(io_toIbuffer_bits_exceptionType_15),
    .io_toIbuffer_bits_crossPageIPFFix_0(io_toIbuffer_bits_crossPageIPFFix_0),
    .io_toIbuffer_bits_crossPageIPFFix_1(io_toIbuffer_bits_crossPageIPFFix_1),
    .io_toIbuffer_bits_crossPageIPFFix_2(io_toIbuffer_bits_crossPageIPFFix_2),
    .io_toIbuffer_bits_crossPageIPFFix_3(io_toIbuffer_bits_crossPageIPFFix_3),
    .io_toIbuffer_bits_crossPageIPFFix_4(io_toIbuffer_bits_crossPageIPFFix_4),
    .io_toIbuffer_bits_crossPageIPFFix_5(io_toIbuffer_bits_crossPageIPFFix_5),
    .io_toIbuffer_bits_crossPageIPFFix_6(io_toIbuffer_bits_crossPageIPFFix_6),
    .io_toIbuffer_bits_crossPageIPFFix_7(io_toIbuffer_bits_crossPageIPFFix_7),
    .io_toIbuffer_bits_crossPageIPFFix_8(io_toIbuffer_bits_crossPageIPFFix_8),
    .io_toIbuffer_bits_crossPageIPFFix_9(io_toIbuffer_bits_crossPageIPFFix_9),
    .io_toIbuffer_bits_crossPageIPFFix_10(io_toIbuffer_bits_crossPageIPFFix_10),
    .io_toIbuffer_bits_crossPageIPFFix_11(io_toIbuffer_bits_crossPageIPFFix_11),
    .io_toIbuffer_bits_crossPageIPFFix_12(io_toIbuffer_bits_crossPageIPFFix_12),
    .io_toIbuffer_bits_crossPageIPFFix_13(io_toIbuffer_bits_crossPageIPFFix_13),
    .io_toIbuffer_bits_crossPageIPFFix_14(io_toIbuffer_bits_crossPageIPFFix_14),
    .io_toIbuffer_bits_crossPageIPFFix_15(io_toIbuffer_bits_crossPageIPFFix_15),
    .io_toIbuffer_bits_illegalInstr_0(io_toIbuffer_bits_illegalInstr_0),
    .io_toIbuffer_bits_illegalInstr_1(io_toIbuffer_bits_illegalInstr_1),
    .io_toIbuffer_bits_illegalInstr_2(io_toIbuffer_bits_illegalInstr_2),
    .io_toIbuffer_bits_illegalInstr_3(io_toIbuffer_bits_illegalInstr_3),
    .io_toIbuffer_bits_illegalInstr_4(io_toIbuffer_bits_illegalInstr_4),
    .io_toIbuffer_bits_illegalInstr_5(io_toIbuffer_bits_illegalInstr_5),
    .io_toIbuffer_bits_illegalInstr_6(io_toIbuffer_bits_illegalInstr_6),
    .io_toIbuffer_bits_illegalInstr_7(io_toIbuffer_bits_illegalInstr_7),
    .io_toIbuffer_bits_illegalInstr_8(io_toIbuffer_bits_illegalInstr_8),
    .io_toIbuffer_bits_illegalInstr_9(io_toIbuffer_bits_illegalInstr_9),
    .io_toIbuffer_bits_illegalInstr_10(io_toIbuffer_bits_illegalInstr_10),
    .io_toIbuffer_bits_illegalInstr_11(io_toIbuffer_bits_illegalInstr_11),
    .io_toIbuffer_bits_illegalInstr_12(io_toIbuffer_bits_illegalInstr_12),
    .io_toIbuffer_bits_illegalInstr_13(io_toIbuffer_bits_illegalInstr_13),
    .io_toIbuffer_bits_illegalInstr_14(io_toIbuffer_bits_illegalInstr_14),
    .io_toIbuffer_bits_illegalInstr_15(io_toIbuffer_bits_illegalInstr_15),
    .io_toIbuffer_bits_triggered_0(io_toIbuffer_bits_triggered_0),
    .io_toIbuffer_bits_triggered_1(io_toIbuffer_bits_triggered_1),
    .io_toIbuffer_bits_triggered_2(io_toIbuffer_bits_triggered_2),
    .io_toIbuffer_bits_triggered_3(io_toIbuffer_bits_triggered_3),
    .io_toIbuffer_bits_triggered_4(io_toIbuffer_bits_triggered_4),
    .io_toIbuffer_bits_triggered_5(io_toIbuffer_bits_triggered_5),
    .io_toIbuffer_bits_triggered_6(io_toIbuffer_bits_triggered_6),
    .io_toIbuffer_bits_triggered_7(io_toIbuffer_bits_triggered_7),
    .io_toIbuffer_bits_triggered_8(io_toIbuffer_bits_triggered_8),
    .io_toIbuffer_bits_triggered_9(io_toIbuffer_bits_triggered_9),
    .io_toIbuffer_bits_triggered_10(io_toIbuffer_bits_triggered_10),
    .io_toIbuffer_bits_triggered_11(io_toIbuffer_bits_triggered_11),
    .io_toIbuffer_bits_triggered_12(io_toIbuffer_bits_triggered_12),
    .io_toIbuffer_bits_triggered_13(io_toIbuffer_bits_triggered_13),
    .io_toIbuffer_bits_triggered_14(io_toIbuffer_bits_triggered_14),
    .io_toIbuffer_bits_triggered_15(io_toIbuffer_bits_triggered_15),
    .io_toIbuffer_bits_isLastInFtqEntry_0(io_toIbuffer_bits_isLastInFtqEntry_0),
    .io_toIbuffer_bits_isLastInFtqEntry_1(io_toIbuffer_bits_isLastInFtqEntry_1),
    .io_toIbuffer_bits_isLastInFtqEntry_2(io_toIbuffer_bits_isLastInFtqEntry_2),
    .io_toIbuffer_bits_isLastInFtqEntry_3(io_toIbuffer_bits_isLastInFtqEntry_3),
    .io_toIbuffer_bits_isLastInFtqEntry_4(io_toIbuffer_bits_isLastInFtqEntry_4),
    .io_toIbuffer_bits_isLastInFtqEntry_5(io_toIbuffer_bits_isLastInFtqEntry_5),
    .io_toIbuffer_bits_isLastInFtqEntry_6(io_toIbuffer_bits_isLastInFtqEntry_6),
    .io_toIbuffer_bits_isLastInFtqEntry_7(io_toIbuffer_bits_isLastInFtqEntry_7),
    .io_toIbuffer_bits_isLastInFtqEntry_8(io_toIbuffer_bits_isLastInFtqEntry_8),
    .io_toIbuffer_bits_isLastInFtqEntry_9(io_toIbuffer_bits_isLastInFtqEntry_9),
    .io_toIbuffer_bits_isLastInFtqEntry_10(io_toIbuffer_bits_isLastInFtqEntry_10),
    .io_toIbuffer_bits_isLastInFtqEntry_11(io_toIbuffer_bits_isLastInFtqEntry_11),
    .io_toIbuffer_bits_isLastInFtqEntry_12(io_toIbuffer_bits_isLastInFtqEntry_12),
    .io_toIbuffer_bits_isLastInFtqEntry_13(io_toIbuffer_bits_isLastInFtqEntry_13),
    .io_toIbuffer_bits_isLastInFtqEntry_14(io_toIbuffer_bits_isLastInFtqEntry_14),
    .io_toIbuffer_bits_isLastInFtqEntry_15(io_toIbuffer_bits_isLastInFtqEntry_15),
    .io_toIbuffer_bits_ftqPtr_flag(io_toIbuffer_bits_ftqPtr_flag),
    .io_toIbuffer_bits_ftqPtr_value(io_toIbuffer_bits_ftqPtr_value),
    .io_toBackend_gpaddrMem_wen(io_toBackend_gpaddrMem_wen),
    .io_toBackend_gpaddrMem_waddr(io_toBackend_gpaddrMem_waddr),
    .io_toBackend_gpaddrMem_wdata_gpaddr(io_toBackend_gpaddrMem_wdata_gpaddr),
    .io_toBackend_gpaddrMem_wdata_isForVSnonLeafPTE(io_toBackend_gpaddrMem_wdata_isForVSnonLeafPTE),
    .io_uncacheInter_fromUncache_valid(io_uncacheInter_fromUncache_valid),
    .io_uncacheInter_fromUncache_bits_data(io_uncacheInter_fromUncache_bits_data),
    .io_uncacheInter_toUncache_ready(io_uncacheInter_toUncache_ready),
    .io_uncacheInter_toUncache_valid(io_uncacheInter_toUncache_valid),
    .io_uncacheInter_toUncache_bits_addr(io_uncacheInter_toUncache_bits_addr),
    .io_frontendTrigger_tUpdate_valid(io_frontendTrigger_tUpdate_valid),
    .io_frontendTrigger_tUpdate_bits_addr(io_frontendTrigger_tUpdate_bits_addr),
    .io_frontendTrigger_tUpdate_bits_tdata_matchType(io_frontendTrigger_tUpdate_bits_tdata_matchType),
    .io_frontendTrigger_tUpdate_bits_tdata_select(io_frontendTrigger_tUpdate_bits_tdata_select),
    .io_frontendTrigger_tUpdate_bits_tdata_action(io_frontendTrigger_tUpdate_bits_tdata_action),
    .io_frontendTrigger_tUpdate_bits_tdata_chain(io_frontendTrigger_tUpdate_bits_tdata_chain),
    .io_frontendTrigger_tUpdate_bits_tdata_tdata2(io_frontendTrigger_tUpdate_bits_tdata_tdata2),
    .io_frontendTrigger_tEnableVec_0(io_frontendTrigger_tEnableVec_0),
    .io_frontendTrigger_tEnableVec_1(io_frontendTrigger_tEnableVec_1),
    .io_frontendTrigger_tEnableVec_2(io_frontendTrigger_tEnableVec_2),
    .io_frontendTrigger_tEnableVec_3(io_frontendTrigger_tEnableVec_3),
    .io_frontendTrigger_debugMode(io_frontendTrigger_debugMode),
    .io_frontendTrigger_triggerCanRaiseBpExp(io_frontendTrigger_triggerCanRaiseBpExp),
    .io_rob_commits_0_valid(io_rob_commits_0_valid),
    .io_rob_commits_0_bits_ftqIdx_flag(io_rob_commits_0_bits_ftqIdx_flag),
    .io_rob_commits_0_bits_ftqIdx_value(io_rob_commits_0_bits_ftqIdx_value),
    .io_rob_commits_0_bits_ftqOffset(io_rob_commits_0_bits_ftqOffset),
    .io_rob_commits_1_valid(io_rob_commits_1_valid),
    .io_rob_commits_1_bits_ftqIdx_flag(io_rob_commits_1_bits_ftqIdx_flag),
    .io_rob_commits_1_bits_ftqIdx_value(io_rob_commits_1_bits_ftqIdx_value),
    .io_rob_commits_1_bits_ftqOffset(io_rob_commits_1_bits_ftqOffset),
    .io_rob_commits_2_valid(io_rob_commits_2_valid),
    .io_rob_commits_2_bits_ftqIdx_flag(io_rob_commits_2_bits_ftqIdx_flag),
    .io_rob_commits_2_bits_ftqIdx_value(io_rob_commits_2_bits_ftqIdx_value),
    .io_rob_commits_2_bits_ftqOffset(io_rob_commits_2_bits_ftqOffset),
    .io_rob_commits_3_valid(io_rob_commits_3_valid),
    .io_rob_commits_3_bits_ftqIdx_flag(io_rob_commits_3_bits_ftqIdx_flag),
    .io_rob_commits_3_bits_ftqIdx_value(io_rob_commits_3_bits_ftqIdx_value),
    .io_rob_commits_3_bits_ftqOffset(io_rob_commits_3_bits_ftqOffset),
    .io_rob_commits_4_valid(io_rob_commits_4_valid),
    .io_rob_commits_4_bits_ftqIdx_flag(io_rob_commits_4_bits_ftqIdx_flag),
    .io_rob_commits_4_bits_ftqIdx_value(io_rob_commits_4_bits_ftqIdx_value),
    .io_rob_commits_4_bits_ftqOffset(io_rob_commits_4_bits_ftqOffset),
    .io_rob_commits_5_valid(io_rob_commits_5_valid),
    .io_rob_commits_5_bits_ftqIdx_flag(io_rob_commits_5_bits_ftqIdx_flag),
    .io_rob_commits_5_bits_ftqIdx_value(io_rob_commits_5_bits_ftqIdx_value),
    .io_rob_commits_5_bits_ftqOffset(io_rob_commits_5_bits_ftqOffset),
    .io_rob_commits_6_valid(io_rob_commits_6_valid),
    .io_rob_commits_6_bits_ftqIdx_flag(io_rob_commits_6_bits_ftqIdx_flag),
    .io_rob_commits_6_bits_ftqIdx_value(io_rob_commits_6_bits_ftqIdx_value),
    .io_rob_commits_6_bits_ftqOffset(io_rob_commits_6_bits_ftqOffset),
    .io_rob_commits_7_valid(io_rob_commits_7_valid),
    .io_rob_commits_7_bits_ftqIdx_flag(io_rob_commits_7_bits_ftqIdx_flag),
    .io_rob_commits_7_bits_ftqIdx_value(io_rob_commits_7_bits_ftqIdx_value),
    .io_rob_commits_7_bits_ftqOffset(io_rob_commits_7_bits_ftqOffset),
    .io_iTLBInter_req_ready(io_iTLBInter_req_ready),
    .io_iTLBInter_req_valid(io_iTLBInter_req_valid),
    .io_iTLBInter_req_bits_vaddr(io_iTLBInter_req_bits_vaddr),
    .io_iTLBInter_resp_ready(io_iTLBInter_resp_ready),
    .io_iTLBInter_resp_valid(io_iTLBInter_resp_valid),
    .io_iTLBInter_resp_bits_paddr_0(io_iTLBInter_resp_bits_paddr_0),
    .io_iTLBInter_resp_bits_gpaddr_0(io_iTLBInter_resp_bits_gpaddr_0),
    .io_iTLBInter_resp_bits_pbmt_0(io_iTLBInter_resp_bits_pbmt_0),
    .io_iTLBInter_resp_bits_isForVSnonLeafPTE(io_iTLBInter_resp_bits_isForVSnonLeafPTE),
    .io_iTLBInter_resp_bits_excp_0_gpf_instr(io_iTLBInter_resp_bits_excp_0_gpf_instr),
    .io_iTLBInter_resp_bits_excp_0_pf_instr(io_iTLBInter_resp_bits_excp_0_pf_instr),
    .io_iTLBInter_resp_bits_excp_0_af_instr(io_iTLBInter_resp_bits_excp_0_af_instr),
    .io_pmp_req_bits_addr(io_pmp_req_bits_addr),
    .io_pmp_resp_instr(io_pmp_resp_instr),
    .io_pmp_resp_mmio(io_pmp_resp_mmio),
    .io_mmioCommitRead_mmioFtqPtr_flag(io_mmioCommitRead_mmioFtqPtr_flag),
    .io_mmioCommitRead_mmioFtqPtr_value(io_mmioCommitRead_mmioFtqPtr_value),
    .io_mmioCommitRead_mmioLastCommit(io_mmioCommitRead_mmioLastCommit),
    .io_csr_fsIsOff(io_csr_fsIsOff),
    .io_perf_0_value(io_perf_0_value),
    .io_perf_1_value(io_perf_1_value),
    .io_perf_2_value(io_perf_2_value),
    .io_perf_3_value(io_perf_3_value),
    .io_perf_4_value(io_perf_4_value),
    .io_perf_5_value(io_perf_5_value),
    .io_perf_6_value(io_perf_6_value),
    .io_perf_7_value(io_perf_7_value),
    .io_perf_8_value(io_perf_8_value),
    .io_perf_9_value(io_perf_9_value),
    .io_perf_10_value(io_perf_10_value),
    .io_perf_11_value(io_perf_11_value),
    .io_perf_12_value(io_perf_12_value)
 );


endmodule

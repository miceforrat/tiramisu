module PredChecker_top;

  logic  clock;
  logic  io_in_ftqOffset_valid;
  logic [3:0] io_in_ftqOffset_bits;
  logic [63:0] io_in_jumpOffset_0;
  logic [63:0] io_in_jumpOffset_1;
  logic [63:0] io_in_jumpOffset_2;
  logic [63:0] io_in_jumpOffset_3;
  logic [63:0] io_in_jumpOffset_4;
  logic [63:0] io_in_jumpOffset_5;
  logic [63:0] io_in_jumpOffset_6;
  logic [63:0] io_in_jumpOffset_7;
  logic [63:0] io_in_jumpOffset_8;
  logic [63:0] io_in_jumpOffset_9;
  logic [63:0] io_in_jumpOffset_10;
  logic [63:0] io_in_jumpOffset_11;
  logic [63:0] io_in_jumpOffset_12;
  logic [63:0] io_in_jumpOffset_13;
  logic [63:0] io_in_jumpOffset_14;
  logic [63:0] io_in_jumpOffset_15;
  logic [49:0] io_in_target;
  logic  io_in_instrRange_0;
  logic  io_in_instrRange_1;
  logic  io_in_instrRange_2;
  logic  io_in_instrRange_3;
  logic  io_in_instrRange_4;
  logic  io_in_instrRange_5;
  logic  io_in_instrRange_6;
  logic  io_in_instrRange_7;
  logic  io_in_instrRange_8;
  logic  io_in_instrRange_9;
  logic  io_in_instrRange_10;
  logic  io_in_instrRange_11;
  logic  io_in_instrRange_12;
  logic  io_in_instrRange_13;
  logic  io_in_instrRange_14;
  logic  io_in_instrRange_15;
  logic  io_in_instrValid_0;
  logic  io_in_instrValid_1;
  logic  io_in_instrValid_2;
  logic  io_in_instrValid_3;
  logic  io_in_instrValid_4;
  logic  io_in_instrValid_5;
  logic  io_in_instrValid_6;
  logic  io_in_instrValid_7;
  logic  io_in_instrValid_8;
  logic  io_in_instrValid_9;
  logic  io_in_instrValid_10;
  logic  io_in_instrValid_11;
  logic  io_in_instrValid_12;
  logic  io_in_instrValid_13;
  logic  io_in_instrValid_14;
  logic  io_in_instrValid_15;
  logic  io_in_pds_0_isRVC;
  logic [1:0] io_in_pds_0_brType;
  logic  io_in_pds_0_isRet;
  logic  io_in_pds_1_isRVC;
  logic [1:0] io_in_pds_1_brType;
  logic  io_in_pds_1_isRet;
  logic  io_in_pds_2_isRVC;
  logic [1:0] io_in_pds_2_brType;
  logic  io_in_pds_2_isRet;
  logic  io_in_pds_3_isRVC;
  logic [1:0] io_in_pds_3_brType;
  logic  io_in_pds_3_isRet;
  logic  io_in_pds_4_isRVC;
  logic [1:0] io_in_pds_4_brType;
  logic  io_in_pds_4_isRet;
  logic  io_in_pds_5_isRVC;
  logic [1:0] io_in_pds_5_brType;
  logic  io_in_pds_5_isRet;
  logic  io_in_pds_6_isRVC;
  logic [1:0] io_in_pds_6_brType;
  logic  io_in_pds_6_isRet;
  logic  io_in_pds_7_isRVC;
  logic [1:0] io_in_pds_7_brType;
  logic  io_in_pds_7_isRet;
  logic  io_in_pds_8_isRVC;
  logic [1:0] io_in_pds_8_brType;
  logic  io_in_pds_8_isRet;
  logic  io_in_pds_9_isRVC;
  logic [1:0] io_in_pds_9_brType;
  logic  io_in_pds_9_isRet;
  logic  io_in_pds_10_isRVC;
  logic [1:0] io_in_pds_10_brType;
  logic  io_in_pds_10_isRet;
  logic  io_in_pds_11_isRVC;
  logic [1:0] io_in_pds_11_brType;
  logic  io_in_pds_11_isRet;
  logic  io_in_pds_12_isRVC;
  logic [1:0] io_in_pds_12_brType;
  logic  io_in_pds_12_isRet;
  logic  io_in_pds_13_isRVC;
  logic [1:0] io_in_pds_13_brType;
  logic  io_in_pds_13_isRet;
  logic  io_in_pds_14_isRVC;
  logic [1:0] io_in_pds_14_brType;
  logic  io_in_pds_14_isRet;
  logic  io_in_pds_15_isRVC;
  logic [1:0] io_in_pds_15_brType;
  logic  io_in_pds_15_isRet;
  logic [49:0] io_in_pc_0;
  logic [49:0] io_in_pc_1;
  logic [49:0] io_in_pc_2;
  logic [49:0] io_in_pc_3;
  logic [49:0] io_in_pc_4;
  logic [49:0] io_in_pc_5;
  logic [49:0] io_in_pc_6;
  logic [49:0] io_in_pc_7;
  logic [49:0] io_in_pc_8;
  logic [49:0] io_in_pc_9;
  logic [49:0] io_in_pc_10;
  logic [49:0] io_in_pc_11;
  logic [49:0] io_in_pc_12;
  logic [49:0] io_in_pc_13;
  logic [49:0] io_in_pc_14;
  logic [49:0] io_in_pc_15;
  logic  io_in_fire_in;
  logic  io_out_stage1Out_fixedRange_0;
  logic  io_out_stage1Out_fixedRange_1;
  logic  io_out_stage1Out_fixedRange_2;
  logic  io_out_stage1Out_fixedRange_3;
  logic  io_out_stage1Out_fixedRange_4;
  logic  io_out_stage1Out_fixedRange_5;
  logic  io_out_stage1Out_fixedRange_6;
  logic  io_out_stage1Out_fixedRange_7;
  logic  io_out_stage1Out_fixedRange_8;
  logic  io_out_stage1Out_fixedRange_9;
  logic  io_out_stage1Out_fixedRange_10;
  logic  io_out_stage1Out_fixedRange_11;
  logic  io_out_stage1Out_fixedRange_12;
  logic  io_out_stage1Out_fixedRange_13;
  logic  io_out_stage1Out_fixedRange_14;
  logic  io_out_stage1Out_fixedRange_15;
  logic  io_out_stage1Out_fixedTaken_0;
  logic  io_out_stage1Out_fixedTaken_1;
  logic  io_out_stage1Out_fixedTaken_2;
  logic  io_out_stage1Out_fixedTaken_3;
  logic  io_out_stage1Out_fixedTaken_4;
  logic  io_out_stage1Out_fixedTaken_5;
  logic  io_out_stage1Out_fixedTaken_6;
  logic  io_out_stage1Out_fixedTaken_7;
  logic  io_out_stage1Out_fixedTaken_8;
  logic  io_out_stage1Out_fixedTaken_9;
  logic  io_out_stage1Out_fixedTaken_10;
  logic  io_out_stage1Out_fixedTaken_11;
  logic  io_out_stage1Out_fixedTaken_12;
  logic  io_out_stage1Out_fixedTaken_13;
  logic  io_out_stage1Out_fixedTaken_14;
  logic  io_out_stage1Out_fixedTaken_15;
  logic [49:0] io_out_stage2Out_fixedTarget_0;
  logic [49:0] io_out_stage2Out_fixedTarget_1;
  logic [49:0] io_out_stage2Out_fixedTarget_2;
  logic [49:0] io_out_stage2Out_fixedTarget_3;
  logic [49:0] io_out_stage2Out_fixedTarget_4;
  logic [49:0] io_out_stage2Out_fixedTarget_5;
  logic [49:0] io_out_stage2Out_fixedTarget_6;
  logic [49:0] io_out_stage2Out_fixedTarget_7;
  logic [49:0] io_out_stage2Out_fixedTarget_8;
  logic [49:0] io_out_stage2Out_fixedTarget_9;
  logic [49:0] io_out_stage2Out_fixedTarget_10;
  logic [49:0] io_out_stage2Out_fixedTarget_11;
  logic [49:0] io_out_stage2Out_fixedTarget_12;
  logic [49:0] io_out_stage2Out_fixedTarget_13;
  logic [49:0] io_out_stage2Out_fixedTarget_14;
  logic [49:0] io_out_stage2Out_fixedTarget_15;
  logic [49:0] io_out_stage2Out_jalTarget_0;
  logic [49:0] io_out_stage2Out_jalTarget_1;
  logic [49:0] io_out_stage2Out_jalTarget_2;
  logic [49:0] io_out_stage2Out_jalTarget_3;
  logic [49:0] io_out_stage2Out_jalTarget_4;
  logic [49:0] io_out_stage2Out_jalTarget_5;
  logic [49:0] io_out_stage2Out_jalTarget_6;
  logic [49:0] io_out_stage2Out_jalTarget_7;
  logic [49:0] io_out_stage2Out_jalTarget_8;
  logic [49:0] io_out_stage2Out_jalTarget_9;
  logic [49:0] io_out_stage2Out_jalTarget_10;
  logic [49:0] io_out_stage2Out_jalTarget_11;
  logic [49:0] io_out_stage2Out_jalTarget_12;
  logic [49:0] io_out_stage2Out_jalTarget_13;
  logic [49:0] io_out_stage2Out_jalTarget_14;
  logic [49:0] io_out_stage2Out_jalTarget_15;
  logic  io_out_stage2Out_fixedMissPred_0;
  logic  io_out_stage2Out_fixedMissPred_1;
  logic  io_out_stage2Out_fixedMissPred_2;
  logic  io_out_stage2Out_fixedMissPred_3;
  logic  io_out_stage2Out_fixedMissPred_4;
  logic  io_out_stage2Out_fixedMissPred_5;
  logic  io_out_stage2Out_fixedMissPred_6;
  logic  io_out_stage2Out_fixedMissPred_7;
  logic  io_out_stage2Out_fixedMissPred_8;
  logic  io_out_stage2Out_fixedMissPred_9;
  logic  io_out_stage2Out_fixedMissPred_10;
  logic  io_out_stage2Out_fixedMissPred_11;
  logic  io_out_stage2Out_fixedMissPred_12;
  logic  io_out_stage2Out_fixedMissPred_13;
  logic  io_out_stage2Out_fixedMissPred_14;
  logic  io_out_stage2Out_fixedMissPred_15;


 PredChecker PredChecker(
    .clock(clock),
    .io_in_ftqOffset_valid(io_in_ftqOffset_valid),
    .io_in_ftqOffset_bits(io_in_ftqOffset_bits),
    .io_in_jumpOffset_0(io_in_jumpOffset_0),
    .io_in_jumpOffset_1(io_in_jumpOffset_1),
    .io_in_jumpOffset_2(io_in_jumpOffset_2),
    .io_in_jumpOffset_3(io_in_jumpOffset_3),
    .io_in_jumpOffset_4(io_in_jumpOffset_4),
    .io_in_jumpOffset_5(io_in_jumpOffset_5),
    .io_in_jumpOffset_6(io_in_jumpOffset_6),
    .io_in_jumpOffset_7(io_in_jumpOffset_7),
    .io_in_jumpOffset_8(io_in_jumpOffset_8),
    .io_in_jumpOffset_9(io_in_jumpOffset_9),
    .io_in_jumpOffset_10(io_in_jumpOffset_10),
    .io_in_jumpOffset_11(io_in_jumpOffset_11),
    .io_in_jumpOffset_12(io_in_jumpOffset_12),
    .io_in_jumpOffset_13(io_in_jumpOffset_13),
    .io_in_jumpOffset_14(io_in_jumpOffset_14),
    .io_in_jumpOffset_15(io_in_jumpOffset_15),
    .io_in_target(io_in_target),
    .io_in_instrRange_0(io_in_instrRange_0),
    .io_in_instrRange_1(io_in_instrRange_1),
    .io_in_instrRange_2(io_in_instrRange_2),
    .io_in_instrRange_3(io_in_instrRange_3),
    .io_in_instrRange_4(io_in_instrRange_4),
    .io_in_instrRange_5(io_in_instrRange_5),
    .io_in_instrRange_6(io_in_instrRange_6),
    .io_in_instrRange_7(io_in_instrRange_7),
    .io_in_instrRange_8(io_in_instrRange_8),
    .io_in_instrRange_9(io_in_instrRange_9),
    .io_in_instrRange_10(io_in_instrRange_10),
    .io_in_instrRange_11(io_in_instrRange_11),
    .io_in_instrRange_12(io_in_instrRange_12),
    .io_in_instrRange_13(io_in_instrRange_13),
    .io_in_instrRange_14(io_in_instrRange_14),
    .io_in_instrRange_15(io_in_instrRange_15),
    .io_in_instrValid_0(io_in_instrValid_0),
    .io_in_instrValid_1(io_in_instrValid_1),
    .io_in_instrValid_2(io_in_instrValid_2),
    .io_in_instrValid_3(io_in_instrValid_3),
    .io_in_instrValid_4(io_in_instrValid_4),
    .io_in_instrValid_5(io_in_instrValid_5),
    .io_in_instrValid_6(io_in_instrValid_6),
    .io_in_instrValid_7(io_in_instrValid_7),
    .io_in_instrValid_8(io_in_instrValid_8),
    .io_in_instrValid_9(io_in_instrValid_9),
    .io_in_instrValid_10(io_in_instrValid_10),
    .io_in_instrValid_11(io_in_instrValid_11),
    .io_in_instrValid_12(io_in_instrValid_12),
    .io_in_instrValid_13(io_in_instrValid_13),
    .io_in_instrValid_14(io_in_instrValid_14),
    .io_in_instrValid_15(io_in_instrValid_15),
    .io_in_pds_0_isRVC(io_in_pds_0_isRVC),
    .io_in_pds_0_brType(io_in_pds_0_brType),
    .io_in_pds_0_isRet(io_in_pds_0_isRet),
    .io_in_pds_1_isRVC(io_in_pds_1_isRVC),
    .io_in_pds_1_brType(io_in_pds_1_brType),
    .io_in_pds_1_isRet(io_in_pds_1_isRet),
    .io_in_pds_2_isRVC(io_in_pds_2_isRVC),
    .io_in_pds_2_brType(io_in_pds_2_brType),
    .io_in_pds_2_isRet(io_in_pds_2_isRet),
    .io_in_pds_3_isRVC(io_in_pds_3_isRVC),
    .io_in_pds_3_brType(io_in_pds_3_brType),
    .io_in_pds_3_isRet(io_in_pds_3_isRet),
    .io_in_pds_4_isRVC(io_in_pds_4_isRVC),
    .io_in_pds_4_brType(io_in_pds_4_brType),
    .io_in_pds_4_isRet(io_in_pds_4_isRet),
    .io_in_pds_5_isRVC(io_in_pds_5_isRVC),
    .io_in_pds_5_brType(io_in_pds_5_brType),
    .io_in_pds_5_isRet(io_in_pds_5_isRet),
    .io_in_pds_6_isRVC(io_in_pds_6_isRVC),
    .io_in_pds_6_brType(io_in_pds_6_brType),
    .io_in_pds_6_isRet(io_in_pds_6_isRet),
    .io_in_pds_7_isRVC(io_in_pds_7_isRVC),
    .io_in_pds_7_brType(io_in_pds_7_brType),
    .io_in_pds_7_isRet(io_in_pds_7_isRet),
    .io_in_pds_8_isRVC(io_in_pds_8_isRVC),
    .io_in_pds_8_brType(io_in_pds_8_brType),
    .io_in_pds_8_isRet(io_in_pds_8_isRet),
    .io_in_pds_9_isRVC(io_in_pds_9_isRVC),
    .io_in_pds_9_brType(io_in_pds_9_brType),
    .io_in_pds_9_isRet(io_in_pds_9_isRet),
    .io_in_pds_10_isRVC(io_in_pds_10_isRVC),
    .io_in_pds_10_brType(io_in_pds_10_brType),
    .io_in_pds_10_isRet(io_in_pds_10_isRet),
    .io_in_pds_11_isRVC(io_in_pds_11_isRVC),
    .io_in_pds_11_brType(io_in_pds_11_brType),
    .io_in_pds_11_isRet(io_in_pds_11_isRet),
    .io_in_pds_12_isRVC(io_in_pds_12_isRVC),
    .io_in_pds_12_brType(io_in_pds_12_brType),
    .io_in_pds_12_isRet(io_in_pds_12_isRet),
    .io_in_pds_13_isRVC(io_in_pds_13_isRVC),
    .io_in_pds_13_brType(io_in_pds_13_brType),
    .io_in_pds_13_isRet(io_in_pds_13_isRet),
    .io_in_pds_14_isRVC(io_in_pds_14_isRVC),
    .io_in_pds_14_brType(io_in_pds_14_brType),
    .io_in_pds_14_isRet(io_in_pds_14_isRet),
    .io_in_pds_15_isRVC(io_in_pds_15_isRVC),
    .io_in_pds_15_brType(io_in_pds_15_brType),
    .io_in_pds_15_isRet(io_in_pds_15_isRet),
    .io_in_pc_0(io_in_pc_0),
    .io_in_pc_1(io_in_pc_1),
    .io_in_pc_2(io_in_pc_2),
    .io_in_pc_3(io_in_pc_3),
    .io_in_pc_4(io_in_pc_4),
    .io_in_pc_5(io_in_pc_5),
    .io_in_pc_6(io_in_pc_6),
    .io_in_pc_7(io_in_pc_7),
    .io_in_pc_8(io_in_pc_8),
    .io_in_pc_9(io_in_pc_9),
    .io_in_pc_10(io_in_pc_10),
    .io_in_pc_11(io_in_pc_11),
    .io_in_pc_12(io_in_pc_12),
    .io_in_pc_13(io_in_pc_13),
    .io_in_pc_14(io_in_pc_14),
    .io_in_pc_15(io_in_pc_15),
    .io_in_fire_in(io_in_fire_in),
    .io_out_stage1Out_fixedRange_0(io_out_stage1Out_fixedRange_0),
    .io_out_stage1Out_fixedRange_1(io_out_stage1Out_fixedRange_1),
    .io_out_stage1Out_fixedRange_2(io_out_stage1Out_fixedRange_2),
    .io_out_stage1Out_fixedRange_3(io_out_stage1Out_fixedRange_3),
    .io_out_stage1Out_fixedRange_4(io_out_stage1Out_fixedRange_4),
    .io_out_stage1Out_fixedRange_5(io_out_stage1Out_fixedRange_5),
    .io_out_stage1Out_fixedRange_6(io_out_stage1Out_fixedRange_6),
    .io_out_stage1Out_fixedRange_7(io_out_stage1Out_fixedRange_7),
    .io_out_stage1Out_fixedRange_8(io_out_stage1Out_fixedRange_8),
    .io_out_stage1Out_fixedRange_9(io_out_stage1Out_fixedRange_9),
    .io_out_stage1Out_fixedRange_10(io_out_stage1Out_fixedRange_10),
    .io_out_stage1Out_fixedRange_11(io_out_stage1Out_fixedRange_11),
    .io_out_stage1Out_fixedRange_12(io_out_stage1Out_fixedRange_12),
    .io_out_stage1Out_fixedRange_13(io_out_stage1Out_fixedRange_13),
    .io_out_stage1Out_fixedRange_14(io_out_stage1Out_fixedRange_14),
    .io_out_stage1Out_fixedRange_15(io_out_stage1Out_fixedRange_15),
    .io_out_stage1Out_fixedTaken_0(io_out_stage1Out_fixedTaken_0),
    .io_out_stage1Out_fixedTaken_1(io_out_stage1Out_fixedTaken_1),
    .io_out_stage1Out_fixedTaken_2(io_out_stage1Out_fixedTaken_2),
    .io_out_stage1Out_fixedTaken_3(io_out_stage1Out_fixedTaken_3),
    .io_out_stage1Out_fixedTaken_4(io_out_stage1Out_fixedTaken_4),
    .io_out_stage1Out_fixedTaken_5(io_out_stage1Out_fixedTaken_5),
    .io_out_stage1Out_fixedTaken_6(io_out_stage1Out_fixedTaken_6),
    .io_out_stage1Out_fixedTaken_7(io_out_stage1Out_fixedTaken_7),
    .io_out_stage1Out_fixedTaken_8(io_out_stage1Out_fixedTaken_8),
    .io_out_stage1Out_fixedTaken_9(io_out_stage1Out_fixedTaken_9),
    .io_out_stage1Out_fixedTaken_10(io_out_stage1Out_fixedTaken_10),
    .io_out_stage1Out_fixedTaken_11(io_out_stage1Out_fixedTaken_11),
    .io_out_stage1Out_fixedTaken_12(io_out_stage1Out_fixedTaken_12),
    .io_out_stage1Out_fixedTaken_13(io_out_stage1Out_fixedTaken_13),
    .io_out_stage1Out_fixedTaken_14(io_out_stage1Out_fixedTaken_14),
    .io_out_stage1Out_fixedTaken_15(io_out_stage1Out_fixedTaken_15),
    .io_out_stage2Out_fixedTarget_0(io_out_stage2Out_fixedTarget_0),
    .io_out_stage2Out_fixedTarget_1(io_out_stage2Out_fixedTarget_1),
    .io_out_stage2Out_fixedTarget_2(io_out_stage2Out_fixedTarget_2),
    .io_out_stage2Out_fixedTarget_3(io_out_stage2Out_fixedTarget_3),
    .io_out_stage2Out_fixedTarget_4(io_out_stage2Out_fixedTarget_4),
    .io_out_stage2Out_fixedTarget_5(io_out_stage2Out_fixedTarget_5),
    .io_out_stage2Out_fixedTarget_6(io_out_stage2Out_fixedTarget_6),
    .io_out_stage2Out_fixedTarget_7(io_out_stage2Out_fixedTarget_7),
    .io_out_stage2Out_fixedTarget_8(io_out_stage2Out_fixedTarget_8),
    .io_out_stage2Out_fixedTarget_9(io_out_stage2Out_fixedTarget_9),
    .io_out_stage2Out_fixedTarget_10(io_out_stage2Out_fixedTarget_10),
    .io_out_stage2Out_fixedTarget_11(io_out_stage2Out_fixedTarget_11),
    .io_out_stage2Out_fixedTarget_12(io_out_stage2Out_fixedTarget_12),
    .io_out_stage2Out_fixedTarget_13(io_out_stage2Out_fixedTarget_13),
    .io_out_stage2Out_fixedTarget_14(io_out_stage2Out_fixedTarget_14),
    .io_out_stage2Out_fixedTarget_15(io_out_stage2Out_fixedTarget_15),
    .io_out_stage2Out_jalTarget_0(io_out_stage2Out_jalTarget_0),
    .io_out_stage2Out_jalTarget_1(io_out_stage2Out_jalTarget_1),
    .io_out_stage2Out_jalTarget_2(io_out_stage2Out_jalTarget_2),
    .io_out_stage2Out_jalTarget_3(io_out_stage2Out_jalTarget_3),
    .io_out_stage2Out_jalTarget_4(io_out_stage2Out_jalTarget_4),
    .io_out_stage2Out_jalTarget_5(io_out_stage2Out_jalTarget_5),
    .io_out_stage2Out_jalTarget_6(io_out_stage2Out_jalTarget_6),
    .io_out_stage2Out_jalTarget_7(io_out_stage2Out_jalTarget_7),
    .io_out_stage2Out_jalTarget_8(io_out_stage2Out_jalTarget_8),
    .io_out_stage2Out_jalTarget_9(io_out_stage2Out_jalTarget_9),
    .io_out_stage2Out_jalTarget_10(io_out_stage2Out_jalTarget_10),
    .io_out_stage2Out_jalTarget_11(io_out_stage2Out_jalTarget_11),
    .io_out_stage2Out_jalTarget_12(io_out_stage2Out_jalTarget_12),
    .io_out_stage2Out_jalTarget_13(io_out_stage2Out_jalTarget_13),
    .io_out_stage2Out_jalTarget_14(io_out_stage2Out_jalTarget_14),
    .io_out_stage2Out_jalTarget_15(io_out_stage2Out_jalTarget_15),
    .io_out_stage2Out_fixedMissPred_0(io_out_stage2Out_fixedMissPred_0),
    .io_out_stage2Out_fixedMissPred_1(io_out_stage2Out_fixedMissPred_1),
    .io_out_stage2Out_fixedMissPred_2(io_out_stage2Out_fixedMissPred_2),
    .io_out_stage2Out_fixedMissPred_3(io_out_stage2Out_fixedMissPred_3),
    .io_out_stage2Out_fixedMissPred_4(io_out_stage2Out_fixedMissPred_4),
    .io_out_stage2Out_fixedMissPred_5(io_out_stage2Out_fixedMissPred_5),
    .io_out_stage2Out_fixedMissPred_6(io_out_stage2Out_fixedMissPred_6),
    .io_out_stage2Out_fixedMissPred_7(io_out_stage2Out_fixedMissPred_7),
    .io_out_stage2Out_fixedMissPred_8(io_out_stage2Out_fixedMissPred_8),
    .io_out_stage2Out_fixedMissPred_9(io_out_stage2Out_fixedMissPred_9),
    .io_out_stage2Out_fixedMissPred_10(io_out_stage2Out_fixedMissPred_10),
    .io_out_stage2Out_fixedMissPred_11(io_out_stage2Out_fixedMissPred_11),
    .io_out_stage2Out_fixedMissPred_12(io_out_stage2Out_fixedMissPred_12),
    .io_out_stage2Out_fixedMissPred_13(io_out_stage2Out_fixedMissPred_13),
    .io_out_stage2Out_fixedMissPred_14(io_out_stage2Out_fixedMissPred_14),
    .io_out_stage2Out_fixedMissPred_15(io_out_stage2Out_fixedMissPred_15)
 );


  export "DPI-C" function get_clockxxPfBDHPCKVf7;
  export "DPI-C" function set_clockxxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_ftqOffset_validxxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_ftqOffset_validxxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_ftqOffset_bitsxxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_ftqOffset_bitsxxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_jumpOffset_0xxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_jumpOffset_0xxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_jumpOffset_1xxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_jumpOffset_1xxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_jumpOffset_2xxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_jumpOffset_2xxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_jumpOffset_3xxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_jumpOffset_3xxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_jumpOffset_4xxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_jumpOffset_4xxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_jumpOffset_5xxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_jumpOffset_5xxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_jumpOffset_6xxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_jumpOffset_6xxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_jumpOffset_7xxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_jumpOffset_7xxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_jumpOffset_8xxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_jumpOffset_8xxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_jumpOffset_9xxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_jumpOffset_9xxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_jumpOffset_10xxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_jumpOffset_10xxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_jumpOffset_11xxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_jumpOffset_11xxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_jumpOffset_12xxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_jumpOffset_12xxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_jumpOffset_13xxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_jumpOffset_13xxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_jumpOffset_14xxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_jumpOffset_14xxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_jumpOffset_15xxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_jumpOffset_15xxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_targetxxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_targetxxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_instrRange_0xxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_instrRange_0xxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_instrRange_1xxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_instrRange_1xxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_instrRange_2xxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_instrRange_2xxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_instrRange_3xxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_instrRange_3xxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_instrRange_4xxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_instrRange_4xxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_instrRange_5xxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_instrRange_5xxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_instrRange_6xxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_instrRange_6xxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_instrRange_7xxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_instrRange_7xxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_instrRange_8xxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_instrRange_8xxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_instrRange_9xxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_instrRange_9xxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_instrRange_10xxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_instrRange_10xxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_instrRange_11xxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_instrRange_11xxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_instrRange_12xxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_instrRange_12xxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_instrRange_13xxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_instrRange_13xxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_instrRange_14xxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_instrRange_14xxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_instrRange_15xxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_instrRange_15xxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_instrValid_0xxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_instrValid_0xxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_instrValid_1xxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_instrValid_1xxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_instrValid_2xxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_instrValid_2xxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_instrValid_3xxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_instrValid_3xxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_instrValid_4xxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_instrValid_4xxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_instrValid_5xxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_instrValid_5xxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_instrValid_6xxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_instrValid_6xxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_instrValid_7xxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_instrValid_7xxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_instrValid_8xxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_instrValid_8xxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_instrValid_9xxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_instrValid_9xxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_instrValid_10xxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_instrValid_10xxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_instrValid_11xxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_instrValid_11xxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_instrValid_12xxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_instrValid_12xxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_instrValid_13xxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_instrValid_13xxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_instrValid_14xxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_instrValid_14xxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_instrValid_15xxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_instrValid_15xxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_pds_0_isRVCxxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_pds_0_isRVCxxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_pds_0_brTypexxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_pds_0_brTypexxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_pds_0_isRetxxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_pds_0_isRetxxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_pds_1_isRVCxxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_pds_1_isRVCxxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_pds_1_brTypexxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_pds_1_brTypexxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_pds_1_isRetxxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_pds_1_isRetxxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_pds_2_isRVCxxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_pds_2_isRVCxxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_pds_2_brTypexxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_pds_2_brTypexxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_pds_2_isRetxxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_pds_2_isRetxxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_pds_3_isRVCxxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_pds_3_isRVCxxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_pds_3_brTypexxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_pds_3_brTypexxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_pds_3_isRetxxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_pds_3_isRetxxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_pds_4_isRVCxxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_pds_4_isRVCxxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_pds_4_brTypexxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_pds_4_brTypexxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_pds_4_isRetxxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_pds_4_isRetxxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_pds_5_isRVCxxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_pds_5_isRVCxxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_pds_5_brTypexxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_pds_5_brTypexxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_pds_5_isRetxxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_pds_5_isRetxxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_pds_6_isRVCxxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_pds_6_isRVCxxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_pds_6_brTypexxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_pds_6_brTypexxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_pds_6_isRetxxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_pds_6_isRetxxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_pds_7_isRVCxxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_pds_7_isRVCxxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_pds_7_brTypexxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_pds_7_brTypexxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_pds_7_isRetxxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_pds_7_isRetxxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_pds_8_isRVCxxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_pds_8_isRVCxxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_pds_8_brTypexxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_pds_8_brTypexxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_pds_8_isRetxxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_pds_8_isRetxxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_pds_9_isRVCxxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_pds_9_isRVCxxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_pds_9_brTypexxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_pds_9_brTypexxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_pds_9_isRetxxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_pds_9_isRetxxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_pds_10_isRVCxxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_pds_10_isRVCxxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_pds_10_brTypexxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_pds_10_brTypexxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_pds_10_isRetxxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_pds_10_isRetxxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_pds_11_isRVCxxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_pds_11_isRVCxxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_pds_11_brTypexxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_pds_11_brTypexxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_pds_11_isRetxxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_pds_11_isRetxxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_pds_12_isRVCxxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_pds_12_isRVCxxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_pds_12_brTypexxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_pds_12_brTypexxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_pds_12_isRetxxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_pds_12_isRetxxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_pds_13_isRVCxxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_pds_13_isRVCxxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_pds_13_brTypexxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_pds_13_brTypexxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_pds_13_isRetxxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_pds_13_isRetxxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_pds_14_isRVCxxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_pds_14_isRVCxxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_pds_14_brTypexxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_pds_14_brTypexxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_pds_14_isRetxxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_pds_14_isRetxxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_pds_15_isRVCxxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_pds_15_isRVCxxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_pds_15_brTypexxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_pds_15_brTypexxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_pds_15_isRetxxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_pds_15_isRetxxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_pc_0xxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_pc_0xxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_pc_1xxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_pc_1xxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_pc_2xxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_pc_2xxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_pc_3xxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_pc_3xxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_pc_4xxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_pc_4xxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_pc_5xxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_pc_5xxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_pc_6xxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_pc_6xxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_pc_7xxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_pc_7xxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_pc_8xxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_pc_8xxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_pc_9xxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_pc_9xxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_pc_10xxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_pc_10xxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_pc_11xxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_pc_11xxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_pc_12xxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_pc_12xxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_pc_13xxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_pc_13xxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_pc_14xxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_pc_14xxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_pc_15xxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_pc_15xxPfBDHPCKVf7;
  export "DPI-C" function get_io_in_fire_inxxPfBDHPCKVf7;
  export "DPI-C" function set_io_in_fire_inxxPfBDHPCKVf7;
  export "DPI-C" function get_io_out_stage1Out_fixedRange_0xxPfBDHPCKVf7;
  export "DPI-C" function set_io_out_stage1Out_fixedRange_0xxPfBDHPCKVf7;
  export "DPI-C" function get_io_out_stage1Out_fixedRange_1xxPfBDHPCKVf7;
  export "DPI-C" function set_io_out_stage1Out_fixedRange_1xxPfBDHPCKVf7;
  export "DPI-C" function get_io_out_stage1Out_fixedRange_2xxPfBDHPCKVf7;
  export "DPI-C" function set_io_out_stage1Out_fixedRange_2xxPfBDHPCKVf7;
  export "DPI-C" function get_io_out_stage1Out_fixedRange_3xxPfBDHPCKVf7;
  export "DPI-C" function set_io_out_stage1Out_fixedRange_3xxPfBDHPCKVf7;
  export "DPI-C" function get_io_out_stage1Out_fixedRange_4xxPfBDHPCKVf7;
  export "DPI-C" function set_io_out_stage1Out_fixedRange_4xxPfBDHPCKVf7;
  export "DPI-C" function get_io_out_stage1Out_fixedRange_5xxPfBDHPCKVf7;
  export "DPI-C" function set_io_out_stage1Out_fixedRange_5xxPfBDHPCKVf7;
  export "DPI-C" function get_io_out_stage1Out_fixedRange_6xxPfBDHPCKVf7;
  export "DPI-C" function set_io_out_stage1Out_fixedRange_6xxPfBDHPCKVf7;
  export "DPI-C" function get_io_out_stage1Out_fixedRange_7xxPfBDHPCKVf7;
  export "DPI-C" function set_io_out_stage1Out_fixedRange_7xxPfBDHPCKVf7;
  export "DPI-C" function get_io_out_stage1Out_fixedRange_8xxPfBDHPCKVf7;
  export "DPI-C" function set_io_out_stage1Out_fixedRange_8xxPfBDHPCKVf7;
  export "DPI-C" function get_io_out_stage1Out_fixedRange_9xxPfBDHPCKVf7;
  export "DPI-C" function set_io_out_stage1Out_fixedRange_9xxPfBDHPCKVf7;
  export "DPI-C" function get_io_out_stage1Out_fixedRange_10xxPfBDHPCKVf7;
  export "DPI-C" function set_io_out_stage1Out_fixedRange_10xxPfBDHPCKVf7;
  export "DPI-C" function get_io_out_stage1Out_fixedRange_11xxPfBDHPCKVf7;
  export "DPI-C" function set_io_out_stage1Out_fixedRange_11xxPfBDHPCKVf7;
  export "DPI-C" function get_io_out_stage1Out_fixedRange_12xxPfBDHPCKVf7;
  export "DPI-C" function set_io_out_stage1Out_fixedRange_12xxPfBDHPCKVf7;
  export "DPI-C" function get_io_out_stage1Out_fixedRange_13xxPfBDHPCKVf7;
  export "DPI-C" function set_io_out_stage1Out_fixedRange_13xxPfBDHPCKVf7;
  export "DPI-C" function get_io_out_stage1Out_fixedRange_14xxPfBDHPCKVf7;
  export "DPI-C" function set_io_out_stage1Out_fixedRange_14xxPfBDHPCKVf7;
  export "DPI-C" function get_io_out_stage1Out_fixedRange_15xxPfBDHPCKVf7;
  export "DPI-C" function set_io_out_stage1Out_fixedRange_15xxPfBDHPCKVf7;
  export "DPI-C" function get_io_out_stage1Out_fixedTaken_0xxPfBDHPCKVf7;
  export "DPI-C" function set_io_out_stage1Out_fixedTaken_0xxPfBDHPCKVf7;
  export "DPI-C" function get_io_out_stage1Out_fixedTaken_1xxPfBDHPCKVf7;
  export "DPI-C" function set_io_out_stage1Out_fixedTaken_1xxPfBDHPCKVf7;
  export "DPI-C" function get_io_out_stage1Out_fixedTaken_2xxPfBDHPCKVf7;
  export "DPI-C" function set_io_out_stage1Out_fixedTaken_2xxPfBDHPCKVf7;
  export "DPI-C" function get_io_out_stage1Out_fixedTaken_3xxPfBDHPCKVf7;
  export "DPI-C" function set_io_out_stage1Out_fixedTaken_3xxPfBDHPCKVf7;
  export "DPI-C" function get_io_out_stage1Out_fixedTaken_4xxPfBDHPCKVf7;
  export "DPI-C" function set_io_out_stage1Out_fixedTaken_4xxPfBDHPCKVf7;
  export "DPI-C" function get_io_out_stage1Out_fixedTaken_5xxPfBDHPCKVf7;
  export "DPI-C" function set_io_out_stage1Out_fixedTaken_5xxPfBDHPCKVf7;
  export "DPI-C" function get_io_out_stage1Out_fixedTaken_6xxPfBDHPCKVf7;
  export "DPI-C" function set_io_out_stage1Out_fixedTaken_6xxPfBDHPCKVf7;
  export "DPI-C" function get_io_out_stage1Out_fixedTaken_7xxPfBDHPCKVf7;
  export "DPI-C" function set_io_out_stage1Out_fixedTaken_7xxPfBDHPCKVf7;
  export "DPI-C" function get_io_out_stage1Out_fixedTaken_8xxPfBDHPCKVf7;
  export "DPI-C" function set_io_out_stage1Out_fixedTaken_8xxPfBDHPCKVf7;
  export "DPI-C" function get_io_out_stage1Out_fixedTaken_9xxPfBDHPCKVf7;
  export "DPI-C" function set_io_out_stage1Out_fixedTaken_9xxPfBDHPCKVf7;
  export "DPI-C" function get_io_out_stage1Out_fixedTaken_10xxPfBDHPCKVf7;
  export "DPI-C" function set_io_out_stage1Out_fixedTaken_10xxPfBDHPCKVf7;
  export "DPI-C" function get_io_out_stage1Out_fixedTaken_11xxPfBDHPCKVf7;
  export "DPI-C" function set_io_out_stage1Out_fixedTaken_11xxPfBDHPCKVf7;
  export "DPI-C" function get_io_out_stage1Out_fixedTaken_12xxPfBDHPCKVf7;
  export "DPI-C" function set_io_out_stage1Out_fixedTaken_12xxPfBDHPCKVf7;
  export "DPI-C" function get_io_out_stage1Out_fixedTaken_13xxPfBDHPCKVf7;
  export "DPI-C" function set_io_out_stage1Out_fixedTaken_13xxPfBDHPCKVf7;
  export "DPI-C" function get_io_out_stage1Out_fixedTaken_14xxPfBDHPCKVf7;
  export "DPI-C" function set_io_out_stage1Out_fixedTaken_14xxPfBDHPCKVf7;
  export "DPI-C" function get_io_out_stage1Out_fixedTaken_15xxPfBDHPCKVf7;
  export "DPI-C" function set_io_out_stage1Out_fixedTaken_15xxPfBDHPCKVf7;
  export "DPI-C" function get_io_out_stage2Out_fixedTarget_0xxPfBDHPCKVf7;
  export "DPI-C" function set_io_out_stage2Out_fixedTarget_0xxPfBDHPCKVf7;
  export "DPI-C" function get_io_out_stage2Out_fixedTarget_1xxPfBDHPCKVf7;
  export "DPI-C" function set_io_out_stage2Out_fixedTarget_1xxPfBDHPCKVf7;
  export "DPI-C" function get_io_out_stage2Out_fixedTarget_2xxPfBDHPCKVf7;
  export "DPI-C" function set_io_out_stage2Out_fixedTarget_2xxPfBDHPCKVf7;
  export "DPI-C" function get_io_out_stage2Out_fixedTarget_3xxPfBDHPCKVf7;
  export "DPI-C" function set_io_out_stage2Out_fixedTarget_3xxPfBDHPCKVf7;
  export "DPI-C" function get_io_out_stage2Out_fixedTarget_4xxPfBDHPCKVf7;
  export "DPI-C" function set_io_out_stage2Out_fixedTarget_4xxPfBDHPCKVf7;
  export "DPI-C" function get_io_out_stage2Out_fixedTarget_5xxPfBDHPCKVf7;
  export "DPI-C" function set_io_out_stage2Out_fixedTarget_5xxPfBDHPCKVf7;
  export "DPI-C" function get_io_out_stage2Out_fixedTarget_6xxPfBDHPCKVf7;
  export "DPI-C" function set_io_out_stage2Out_fixedTarget_6xxPfBDHPCKVf7;
  export "DPI-C" function get_io_out_stage2Out_fixedTarget_7xxPfBDHPCKVf7;
  export "DPI-C" function set_io_out_stage2Out_fixedTarget_7xxPfBDHPCKVf7;
  export "DPI-C" function get_io_out_stage2Out_fixedTarget_8xxPfBDHPCKVf7;
  export "DPI-C" function set_io_out_stage2Out_fixedTarget_8xxPfBDHPCKVf7;
  export "DPI-C" function get_io_out_stage2Out_fixedTarget_9xxPfBDHPCKVf7;
  export "DPI-C" function set_io_out_stage2Out_fixedTarget_9xxPfBDHPCKVf7;
  export "DPI-C" function get_io_out_stage2Out_fixedTarget_10xxPfBDHPCKVf7;
  export "DPI-C" function set_io_out_stage2Out_fixedTarget_10xxPfBDHPCKVf7;
  export "DPI-C" function get_io_out_stage2Out_fixedTarget_11xxPfBDHPCKVf7;
  export "DPI-C" function set_io_out_stage2Out_fixedTarget_11xxPfBDHPCKVf7;
  export "DPI-C" function get_io_out_stage2Out_fixedTarget_12xxPfBDHPCKVf7;
  export "DPI-C" function set_io_out_stage2Out_fixedTarget_12xxPfBDHPCKVf7;
  export "DPI-C" function get_io_out_stage2Out_fixedTarget_13xxPfBDHPCKVf7;
  export "DPI-C" function set_io_out_stage2Out_fixedTarget_13xxPfBDHPCKVf7;
  export "DPI-C" function get_io_out_stage2Out_fixedTarget_14xxPfBDHPCKVf7;
  export "DPI-C" function set_io_out_stage2Out_fixedTarget_14xxPfBDHPCKVf7;
  export "DPI-C" function get_io_out_stage2Out_fixedTarget_15xxPfBDHPCKVf7;
  export "DPI-C" function set_io_out_stage2Out_fixedTarget_15xxPfBDHPCKVf7;
  export "DPI-C" function get_io_out_stage2Out_jalTarget_0xxPfBDHPCKVf7;
  export "DPI-C" function set_io_out_stage2Out_jalTarget_0xxPfBDHPCKVf7;
  export "DPI-C" function get_io_out_stage2Out_jalTarget_1xxPfBDHPCKVf7;
  export "DPI-C" function set_io_out_stage2Out_jalTarget_1xxPfBDHPCKVf7;
  export "DPI-C" function get_io_out_stage2Out_jalTarget_2xxPfBDHPCKVf7;
  export "DPI-C" function set_io_out_stage2Out_jalTarget_2xxPfBDHPCKVf7;
  export "DPI-C" function get_io_out_stage2Out_jalTarget_3xxPfBDHPCKVf7;
  export "DPI-C" function set_io_out_stage2Out_jalTarget_3xxPfBDHPCKVf7;
  export "DPI-C" function get_io_out_stage2Out_jalTarget_4xxPfBDHPCKVf7;
  export "DPI-C" function set_io_out_stage2Out_jalTarget_4xxPfBDHPCKVf7;
  export "DPI-C" function get_io_out_stage2Out_jalTarget_5xxPfBDHPCKVf7;
  export "DPI-C" function set_io_out_stage2Out_jalTarget_5xxPfBDHPCKVf7;
  export "DPI-C" function get_io_out_stage2Out_jalTarget_6xxPfBDHPCKVf7;
  export "DPI-C" function set_io_out_stage2Out_jalTarget_6xxPfBDHPCKVf7;
  export "DPI-C" function get_io_out_stage2Out_jalTarget_7xxPfBDHPCKVf7;
  export "DPI-C" function set_io_out_stage2Out_jalTarget_7xxPfBDHPCKVf7;
  export "DPI-C" function get_io_out_stage2Out_jalTarget_8xxPfBDHPCKVf7;
  export "DPI-C" function set_io_out_stage2Out_jalTarget_8xxPfBDHPCKVf7;
  export "DPI-C" function get_io_out_stage2Out_jalTarget_9xxPfBDHPCKVf7;
  export "DPI-C" function set_io_out_stage2Out_jalTarget_9xxPfBDHPCKVf7;
  export "DPI-C" function get_io_out_stage2Out_jalTarget_10xxPfBDHPCKVf7;
  export "DPI-C" function set_io_out_stage2Out_jalTarget_10xxPfBDHPCKVf7;
  export "DPI-C" function get_io_out_stage2Out_jalTarget_11xxPfBDHPCKVf7;
  export "DPI-C" function set_io_out_stage2Out_jalTarget_11xxPfBDHPCKVf7;
  export "DPI-C" function get_io_out_stage2Out_jalTarget_12xxPfBDHPCKVf7;
  export "DPI-C" function set_io_out_stage2Out_jalTarget_12xxPfBDHPCKVf7;
  export "DPI-C" function get_io_out_stage2Out_jalTarget_13xxPfBDHPCKVf7;
  export "DPI-C" function set_io_out_stage2Out_jalTarget_13xxPfBDHPCKVf7;
  export "DPI-C" function get_io_out_stage2Out_jalTarget_14xxPfBDHPCKVf7;
  export "DPI-C" function set_io_out_stage2Out_jalTarget_14xxPfBDHPCKVf7;
  export "DPI-C" function get_io_out_stage2Out_jalTarget_15xxPfBDHPCKVf7;
  export "DPI-C" function set_io_out_stage2Out_jalTarget_15xxPfBDHPCKVf7;
  export "DPI-C" function get_io_out_stage2Out_fixedMissPred_0xxPfBDHPCKVf7;
  export "DPI-C" function set_io_out_stage2Out_fixedMissPred_0xxPfBDHPCKVf7;
  export "DPI-C" function get_io_out_stage2Out_fixedMissPred_1xxPfBDHPCKVf7;
  export "DPI-C" function set_io_out_stage2Out_fixedMissPred_1xxPfBDHPCKVf7;
  export "DPI-C" function get_io_out_stage2Out_fixedMissPred_2xxPfBDHPCKVf7;
  export "DPI-C" function set_io_out_stage2Out_fixedMissPred_2xxPfBDHPCKVf7;
  export "DPI-C" function get_io_out_stage2Out_fixedMissPred_3xxPfBDHPCKVf7;
  export "DPI-C" function set_io_out_stage2Out_fixedMissPred_3xxPfBDHPCKVf7;
  export "DPI-C" function get_io_out_stage2Out_fixedMissPred_4xxPfBDHPCKVf7;
  export "DPI-C" function set_io_out_stage2Out_fixedMissPred_4xxPfBDHPCKVf7;
  export "DPI-C" function get_io_out_stage2Out_fixedMissPred_5xxPfBDHPCKVf7;
  export "DPI-C" function set_io_out_stage2Out_fixedMissPred_5xxPfBDHPCKVf7;
  export "DPI-C" function get_io_out_stage2Out_fixedMissPred_6xxPfBDHPCKVf7;
  export "DPI-C" function set_io_out_stage2Out_fixedMissPred_6xxPfBDHPCKVf7;
  export "DPI-C" function get_io_out_stage2Out_fixedMissPred_7xxPfBDHPCKVf7;
  export "DPI-C" function set_io_out_stage2Out_fixedMissPred_7xxPfBDHPCKVf7;
  export "DPI-C" function get_io_out_stage2Out_fixedMissPred_8xxPfBDHPCKVf7;
  export "DPI-C" function set_io_out_stage2Out_fixedMissPred_8xxPfBDHPCKVf7;
  export "DPI-C" function get_io_out_stage2Out_fixedMissPred_9xxPfBDHPCKVf7;
  export "DPI-C" function set_io_out_stage2Out_fixedMissPred_9xxPfBDHPCKVf7;
  export "DPI-C" function get_io_out_stage2Out_fixedMissPred_10xxPfBDHPCKVf7;
  export "DPI-C" function set_io_out_stage2Out_fixedMissPred_10xxPfBDHPCKVf7;
  export "DPI-C" function get_io_out_stage2Out_fixedMissPred_11xxPfBDHPCKVf7;
  export "DPI-C" function set_io_out_stage2Out_fixedMissPred_11xxPfBDHPCKVf7;
  export "DPI-C" function get_io_out_stage2Out_fixedMissPred_12xxPfBDHPCKVf7;
  export "DPI-C" function set_io_out_stage2Out_fixedMissPred_12xxPfBDHPCKVf7;
  export "DPI-C" function get_io_out_stage2Out_fixedMissPred_13xxPfBDHPCKVf7;
  export "DPI-C" function set_io_out_stage2Out_fixedMissPred_13xxPfBDHPCKVf7;
  export "DPI-C" function get_io_out_stage2Out_fixedMissPred_14xxPfBDHPCKVf7;
  export "DPI-C" function set_io_out_stage2Out_fixedMissPred_14xxPfBDHPCKVf7;
  export "DPI-C" function get_io_out_stage2Out_fixedMissPred_15xxPfBDHPCKVf7;
  export "DPI-C" function set_io_out_stage2Out_fixedMissPred_15xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_jalFaultVec_0xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_jalFaultVec_1xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_jalFaultVec_2xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_jalFaultVec_3xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_jalFaultVec_4xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_jalFaultVec_5xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_jalFaultVec_6xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_jalFaultVec_7xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_jalFaultVec_8xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_jalFaultVec_9xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_jalFaultVec_10xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_jalFaultVec_11xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_jalFaultVec_12xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_jalFaultVec_13xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_jalFaultVec_14xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_jalFaultVec_15xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_retFaultVec_0xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_retFaultVec_1xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_retFaultVec_2xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_retFaultVec_3xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_retFaultVec_4xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_retFaultVec_5xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_retFaultVec_6xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_retFaultVec_7xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_retFaultVec_8xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_retFaultVec_9xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_retFaultVec_10xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_retFaultVec_11xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_retFaultVec_12xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_retFaultVec_13xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_retFaultVec_14xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_retFaultVec_15xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_remaskFault_0xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_remaskFault_1xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_remaskFault_2xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_remaskFault_3xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_remaskFault_4xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_remaskFault_5xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_remaskFault_6xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_remaskFault_7xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_remaskFault_8xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_remaskFault_9xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_remaskFault_10xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_remaskFault_11xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_remaskFault_12xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_remaskFault_13xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_remaskFault_14xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_fixedRangexxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_fixedRangeNextxxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_instrValidNext_0xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_instrValidNext_1xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_instrValidNext_2xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_instrValidNext_3xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_instrValidNext_4xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_instrValidNext_5xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_instrValidNext_6xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_instrValidNext_7xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_instrValidNext_8xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_instrValidNext_9xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_instrValidNext_10xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_instrValidNext_11xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_instrValidNext_12xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_instrValidNext_13xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_instrValidNext_14xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_instrValidNext_15xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_takenIdxNextxxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_predTakenNextxxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_predTargetNextxxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_jumpTargetsNext_0xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_jumpTargetsNext_1xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_jumpTargetsNext_2xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_jumpTargetsNext_3xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_jumpTargetsNext_4xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_jumpTargetsNext_5xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_jumpTargetsNext_6xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_jumpTargetsNext_7xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_jumpTargetsNext_8xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_jumpTargetsNext_9xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_jumpTargetsNext_10xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_jumpTargetsNext_11xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_jumpTargetsNext_12xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_jumpTargetsNext_13xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_jumpTargetsNext_14xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_jumpTargetsNext_15xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_seqTargetsNext_0xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_seqTargetsNext_1xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_seqTargetsNext_2xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_seqTargetsNext_3xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_seqTargetsNext_4xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_seqTargetsNext_5xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_seqTargetsNext_6xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_seqTargetsNext_7xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_seqTargetsNext_8xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_seqTargetsNext_9xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_seqTargetsNext_10xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_seqTargetsNext_11xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_seqTargetsNext_12xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_seqTargetsNext_13xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_seqTargetsNext_14xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_seqTargetsNext_15xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_pdsNext_0_brTypexxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_pdsNext_1_brTypexxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_pdsNext_2_brTypexxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_pdsNext_3_brTypexxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_pdsNext_4_brTypexxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_pdsNext_5_brTypexxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_pdsNext_6_brTypexxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_pdsNext_7_brTypexxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_pdsNext_8_brTypexxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_pdsNext_9_brTypexxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_pdsNext_10_brTypexxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_pdsNext_11_brTypexxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_pdsNext_12_brTypexxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_pdsNext_13_brTypexxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_pdsNext_14_brTypexxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_pdsNext_15_brTypexxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_jalFaultVecNext_0xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_jalFaultVecNext_1xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_jalFaultVecNext_2xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_jalFaultVecNext_3xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_jalFaultVecNext_4xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_jalFaultVecNext_5xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_jalFaultVecNext_6xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_jalFaultVecNext_7xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_jalFaultVecNext_8xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_jalFaultVecNext_9xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_jalFaultVecNext_10xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_jalFaultVecNext_11xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_jalFaultVecNext_12xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_jalFaultVecNext_13xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_jalFaultVecNext_14xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_jalFaultVecNext_15xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_retFaultVecNext_0xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_retFaultVecNext_1xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_retFaultVecNext_2xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_retFaultVecNext_3xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_retFaultVecNext_4xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_retFaultVecNext_5xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_retFaultVecNext_6xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_retFaultVecNext_7xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_retFaultVecNext_8xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_retFaultVecNext_9xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_retFaultVecNext_10xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_retFaultVecNext_11xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_retFaultVecNext_12xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_retFaultVecNext_13xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_retFaultVecNext_14xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_retFaultVecNext_15xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_notCFITakenNext_0xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_notCFITakenNext_1xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_notCFITakenNext_2xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_notCFITakenNext_3xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_notCFITakenNext_4xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_notCFITakenNext_5xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_notCFITakenNext_6xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_notCFITakenNext_7xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_notCFITakenNext_8xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_notCFITakenNext_9xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_notCFITakenNext_10xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_notCFITakenNext_11xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_notCFITakenNext_12xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_notCFITakenNext_13xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_notCFITakenNext_14xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_notCFITakenNext_15xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_invalidTakenNext_0xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_invalidTakenNext_1xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_invalidTakenNext_2xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_invalidTakenNext_3xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_invalidTakenNext_4xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_invalidTakenNext_5xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_invalidTakenNext_6xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_invalidTakenNext_7xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_invalidTakenNext_8xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_invalidTakenNext_9xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_invalidTakenNext_10xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_invalidTakenNext_11xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_invalidTakenNext_12xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_invalidTakenNext_13xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_invalidTakenNext_14xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_invalidTakenNext_15xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_targetFault_0xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_targetFault_1xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_targetFault_2xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_targetFault_3xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_targetFault_4xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_targetFault_5xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_targetFault_6xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_targetFault_7xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_targetFault_8xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_targetFault_9xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_targetFault_10xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_targetFault_11xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_targetFault_12xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_targetFault_13xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_targetFault_14xxPfBDHPCKVf7;
  export "DPI-C" function get_PredChecker_targetFault_15xxPfBDHPCKVf7;


  function void get_clockxxPfBDHPCKVf7;
    output logic  value;
    value=clock;
  endfunction

  function void set_clockxxPfBDHPCKVf7;
    input logic  value;
    clock=value;
  endfunction

  function void get_io_in_ftqOffset_validxxPfBDHPCKVf7;
    output logic  value;
    value=io_in_ftqOffset_valid;
  endfunction

  function void set_io_in_ftqOffset_validxxPfBDHPCKVf7;
    input logic  value;
    io_in_ftqOffset_valid=value;
  endfunction

  function void get_io_in_ftqOffset_bitsxxPfBDHPCKVf7;
    output logic [3:0] value;
    value=io_in_ftqOffset_bits;
  endfunction

  function void set_io_in_ftqOffset_bitsxxPfBDHPCKVf7;
    input logic [3:0] value;
    io_in_ftqOffset_bits=value;
  endfunction

  function void get_io_in_jumpOffset_0xxPfBDHPCKVf7;
    output logic [63:0] value;
    value=io_in_jumpOffset_0;
  endfunction

  function void set_io_in_jumpOffset_0xxPfBDHPCKVf7;
    input logic [63:0] value;
    io_in_jumpOffset_0=value;
  endfunction

  function void get_io_in_jumpOffset_1xxPfBDHPCKVf7;
    output logic [63:0] value;
    value=io_in_jumpOffset_1;
  endfunction

  function void set_io_in_jumpOffset_1xxPfBDHPCKVf7;
    input logic [63:0] value;
    io_in_jumpOffset_1=value;
  endfunction

  function void get_io_in_jumpOffset_2xxPfBDHPCKVf7;
    output logic [63:0] value;
    value=io_in_jumpOffset_2;
  endfunction

  function void set_io_in_jumpOffset_2xxPfBDHPCKVf7;
    input logic [63:0] value;
    io_in_jumpOffset_2=value;
  endfunction

  function void get_io_in_jumpOffset_3xxPfBDHPCKVf7;
    output logic [63:0] value;
    value=io_in_jumpOffset_3;
  endfunction

  function void set_io_in_jumpOffset_3xxPfBDHPCKVf7;
    input logic [63:0] value;
    io_in_jumpOffset_3=value;
  endfunction

  function void get_io_in_jumpOffset_4xxPfBDHPCKVf7;
    output logic [63:0] value;
    value=io_in_jumpOffset_4;
  endfunction

  function void set_io_in_jumpOffset_4xxPfBDHPCKVf7;
    input logic [63:0] value;
    io_in_jumpOffset_4=value;
  endfunction

  function void get_io_in_jumpOffset_5xxPfBDHPCKVf7;
    output logic [63:0] value;
    value=io_in_jumpOffset_5;
  endfunction

  function void set_io_in_jumpOffset_5xxPfBDHPCKVf7;
    input logic [63:0] value;
    io_in_jumpOffset_5=value;
  endfunction

  function void get_io_in_jumpOffset_6xxPfBDHPCKVf7;
    output logic [63:0] value;
    value=io_in_jumpOffset_6;
  endfunction

  function void set_io_in_jumpOffset_6xxPfBDHPCKVf7;
    input logic [63:0] value;
    io_in_jumpOffset_6=value;
  endfunction

  function void get_io_in_jumpOffset_7xxPfBDHPCKVf7;
    output logic [63:0] value;
    value=io_in_jumpOffset_7;
  endfunction

  function void set_io_in_jumpOffset_7xxPfBDHPCKVf7;
    input logic [63:0] value;
    io_in_jumpOffset_7=value;
  endfunction

  function void get_io_in_jumpOffset_8xxPfBDHPCKVf7;
    output logic [63:0] value;
    value=io_in_jumpOffset_8;
  endfunction

  function void set_io_in_jumpOffset_8xxPfBDHPCKVf7;
    input logic [63:0] value;
    io_in_jumpOffset_8=value;
  endfunction

  function void get_io_in_jumpOffset_9xxPfBDHPCKVf7;
    output logic [63:0] value;
    value=io_in_jumpOffset_9;
  endfunction

  function void set_io_in_jumpOffset_9xxPfBDHPCKVf7;
    input logic [63:0] value;
    io_in_jumpOffset_9=value;
  endfunction

  function void get_io_in_jumpOffset_10xxPfBDHPCKVf7;
    output logic [63:0] value;
    value=io_in_jumpOffset_10;
  endfunction

  function void set_io_in_jumpOffset_10xxPfBDHPCKVf7;
    input logic [63:0] value;
    io_in_jumpOffset_10=value;
  endfunction

  function void get_io_in_jumpOffset_11xxPfBDHPCKVf7;
    output logic [63:0] value;
    value=io_in_jumpOffset_11;
  endfunction

  function void set_io_in_jumpOffset_11xxPfBDHPCKVf7;
    input logic [63:0] value;
    io_in_jumpOffset_11=value;
  endfunction

  function void get_io_in_jumpOffset_12xxPfBDHPCKVf7;
    output logic [63:0] value;
    value=io_in_jumpOffset_12;
  endfunction

  function void set_io_in_jumpOffset_12xxPfBDHPCKVf7;
    input logic [63:0] value;
    io_in_jumpOffset_12=value;
  endfunction

  function void get_io_in_jumpOffset_13xxPfBDHPCKVf7;
    output logic [63:0] value;
    value=io_in_jumpOffset_13;
  endfunction

  function void set_io_in_jumpOffset_13xxPfBDHPCKVf7;
    input logic [63:0] value;
    io_in_jumpOffset_13=value;
  endfunction

  function void get_io_in_jumpOffset_14xxPfBDHPCKVf7;
    output logic [63:0] value;
    value=io_in_jumpOffset_14;
  endfunction

  function void set_io_in_jumpOffset_14xxPfBDHPCKVf7;
    input logic [63:0] value;
    io_in_jumpOffset_14=value;
  endfunction

  function void get_io_in_jumpOffset_15xxPfBDHPCKVf7;
    output logic [63:0] value;
    value=io_in_jumpOffset_15;
  endfunction

  function void set_io_in_jumpOffset_15xxPfBDHPCKVf7;
    input logic [63:0] value;
    io_in_jumpOffset_15=value;
  endfunction

  function void get_io_in_targetxxPfBDHPCKVf7;
    output logic [49:0] value;
    value=io_in_target;
  endfunction

  function void set_io_in_targetxxPfBDHPCKVf7;
    input logic [49:0] value;
    io_in_target=value;
  endfunction

  function void get_io_in_instrRange_0xxPfBDHPCKVf7;
    output logic  value;
    value=io_in_instrRange_0;
  endfunction

  function void set_io_in_instrRange_0xxPfBDHPCKVf7;
    input logic  value;
    io_in_instrRange_0=value;
  endfunction

  function void get_io_in_instrRange_1xxPfBDHPCKVf7;
    output logic  value;
    value=io_in_instrRange_1;
  endfunction

  function void set_io_in_instrRange_1xxPfBDHPCKVf7;
    input logic  value;
    io_in_instrRange_1=value;
  endfunction

  function void get_io_in_instrRange_2xxPfBDHPCKVf7;
    output logic  value;
    value=io_in_instrRange_2;
  endfunction

  function void set_io_in_instrRange_2xxPfBDHPCKVf7;
    input logic  value;
    io_in_instrRange_2=value;
  endfunction

  function void get_io_in_instrRange_3xxPfBDHPCKVf7;
    output logic  value;
    value=io_in_instrRange_3;
  endfunction

  function void set_io_in_instrRange_3xxPfBDHPCKVf7;
    input logic  value;
    io_in_instrRange_3=value;
  endfunction

  function void get_io_in_instrRange_4xxPfBDHPCKVf7;
    output logic  value;
    value=io_in_instrRange_4;
  endfunction

  function void set_io_in_instrRange_4xxPfBDHPCKVf7;
    input logic  value;
    io_in_instrRange_4=value;
  endfunction

  function void get_io_in_instrRange_5xxPfBDHPCKVf7;
    output logic  value;
    value=io_in_instrRange_5;
  endfunction

  function void set_io_in_instrRange_5xxPfBDHPCKVf7;
    input logic  value;
    io_in_instrRange_5=value;
  endfunction

  function void get_io_in_instrRange_6xxPfBDHPCKVf7;
    output logic  value;
    value=io_in_instrRange_6;
  endfunction

  function void set_io_in_instrRange_6xxPfBDHPCKVf7;
    input logic  value;
    io_in_instrRange_6=value;
  endfunction

  function void get_io_in_instrRange_7xxPfBDHPCKVf7;
    output logic  value;
    value=io_in_instrRange_7;
  endfunction

  function void set_io_in_instrRange_7xxPfBDHPCKVf7;
    input logic  value;
    io_in_instrRange_7=value;
  endfunction

  function void get_io_in_instrRange_8xxPfBDHPCKVf7;
    output logic  value;
    value=io_in_instrRange_8;
  endfunction

  function void set_io_in_instrRange_8xxPfBDHPCKVf7;
    input logic  value;
    io_in_instrRange_8=value;
  endfunction

  function void get_io_in_instrRange_9xxPfBDHPCKVf7;
    output logic  value;
    value=io_in_instrRange_9;
  endfunction

  function void set_io_in_instrRange_9xxPfBDHPCKVf7;
    input logic  value;
    io_in_instrRange_9=value;
  endfunction

  function void get_io_in_instrRange_10xxPfBDHPCKVf7;
    output logic  value;
    value=io_in_instrRange_10;
  endfunction

  function void set_io_in_instrRange_10xxPfBDHPCKVf7;
    input logic  value;
    io_in_instrRange_10=value;
  endfunction

  function void get_io_in_instrRange_11xxPfBDHPCKVf7;
    output logic  value;
    value=io_in_instrRange_11;
  endfunction

  function void set_io_in_instrRange_11xxPfBDHPCKVf7;
    input logic  value;
    io_in_instrRange_11=value;
  endfunction

  function void get_io_in_instrRange_12xxPfBDHPCKVf7;
    output logic  value;
    value=io_in_instrRange_12;
  endfunction

  function void set_io_in_instrRange_12xxPfBDHPCKVf7;
    input logic  value;
    io_in_instrRange_12=value;
  endfunction

  function void get_io_in_instrRange_13xxPfBDHPCKVf7;
    output logic  value;
    value=io_in_instrRange_13;
  endfunction

  function void set_io_in_instrRange_13xxPfBDHPCKVf7;
    input logic  value;
    io_in_instrRange_13=value;
  endfunction

  function void get_io_in_instrRange_14xxPfBDHPCKVf7;
    output logic  value;
    value=io_in_instrRange_14;
  endfunction

  function void set_io_in_instrRange_14xxPfBDHPCKVf7;
    input logic  value;
    io_in_instrRange_14=value;
  endfunction

  function void get_io_in_instrRange_15xxPfBDHPCKVf7;
    output logic  value;
    value=io_in_instrRange_15;
  endfunction

  function void set_io_in_instrRange_15xxPfBDHPCKVf7;
    input logic  value;
    io_in_instrRange_15=value;
  endfunction

  function void get_io_in_instrValid_0xxPfBDHPCKVf7;
    output logic  value;
    value=io_in_instrValid_0;
  endfunction

  function void set_io_in_instrValid_0xxPfBDHPCKVf7;
    input logic  value;
    io_in_instrValid_0=value;
  endfunction

  function void get_io_in_instrValid_1xxPfBDHPCKVf7;
    output logic  value;
    value=io_in_instrValid_1;
  endfunction

  function void set_io_in_instrValid_1xxPfBDHPCKVf7;
    input logic  value;
    io_in_instrValid_1=value;
  endfunction

  function void get_io_in_instrValid_2xxPfBDHPCKVf7;
    output logic  value;
    value=io_in_instrValid_2;
  endfunction

  function void set_io_in_instrValid_2xxPfBDHPCKVf7;
    input logic  value;
    io_in_instrValid_2=value;
  endfunction

  function void get_io_in_instrValid_3xxPfBDHPCKVf7;
    output logic  value;
    value=io_in_instrValid_3;
  endfunction

  function void set_io_in_instrValid_3xxPfBDHPCKVf7;
    input logic  value;
    io_in_instrValid_3=value;
  endfunction

  function void get_io_in_instrValid_4xxPfBDHPCKVf7;
    output logic  value;
    value=io_in_instrValid_4;
  endfunction

  function void set_io_in_instrValid_4xxPfBDHPCKVf7;
    input logic  value;
    io_in_instrValid_4=value;
  endfunction

  function void get_io_in_instrValid_5xxPfBDHPCKVf7;
    output logic  value;
    value=io_in_instrValid_5;
  endfunction

  function void set_io_in_instrValid_5xxPfBDHPCKVf7;
    input logic  value;
    io_in_instrValid_5=value;
  endfunction

  function void get_io_in_instrValid_6xxPfBDHPCKVf7;
    output logic  value;
    value=io_in_instrValid_6;
  endfunction

  function void set_io_in_instrValid_6xxPfBDHPCKVf7;
    input logic  value;
    io_in_instrValid_6=value;
  endfunction

  function void get_io_in_instrValid_7xxPfBDHPCKVf7;
    output logic  value;
    value=io_in_instrValid_7;
  endfunction

  function void set_io_in_instrValid_7xxPfBDHPCKVf7;
    input logic  value;
    io_in_instrValid_7=value;
  endfunction

  function void get_io_in_instrValid_8xxPfBDHPCKVf7;
    output logic  value;
    value=io_in_instrValid_8;
  endfunction

  function void set_io_in_instrValid_8xxPfBDHPCKVf7;
    input logic  value;
    io_in_instrValid_8=value;
  endfunction

  function void get_io_in_instrValid_9xxPfBDHPCKVf7;
    output logic  value;
    value=io_in_instrValid_9;
  endfunction

  function void set_io_in_instrValid_9xxPfBDHPCKVf7;
    input logic  value;
    io_in_instrValid_9=value;
  endfunction

  function void get_io_in_instrValid_10xxPfBDHPCKVf7;
    output logic  value;
    value=io_in_instrValid_10;
  endfunction

  function void set_io_in_instrValid_10xxPfBDHPCKVf7;
    input logic  value;
    io_in_instrValid_10=value;
  endfunction

  function void get_io_in_instrValid_11xxPfBDHPCKVf7;
    output logic  value;
    value=io_in_instrValid_11;
  endfunction

  function void set_io_in_instrValid_11xxPfBDHPCKVf7;
    input logic  value;
    io_in_instrValid_11=value;
  endfunction

  function void get_io_in_instrValid_12xxPfBDHPCKVf7;
    output logic  value;
    value=io_in_instrValid_12;
  endfunction

  function void set_io_in_instrValid_12xxPfBDHPCKVf7;
    input logic  value;
    io_in_instrValid_12=value;
  endfunction

  function void get_io_in_instrValid_13xxPfBDHPCKVf7;
    output logic  value;
    value=io_in_instrValid_13;
  endfunction

  function void set_io_in_instrValid_13xxPfBDHPCKVf7;
    input logic  value;
    io_in_instrValid_13=value;
  endfunction

  function void get_io_in_instrValid_14xxPfBDHPCKVf7;
    output logic  value;
    value=io_in_instrValid_14;
  endfunction

  function void set_io_in_instrValid_14xxPfBDHPCKVf7;
    input logic  value;
    io_in_instrValid_14=value;
  endfunction

  function void get_io_in_instrValid_15xxPfBDHPCKVf7;
    output logic  value;
    value=io_in_instrValid_15;
  endfunction

  function void set_io_in_instrValid_15xxPfBDHPCKVf7;
    input logic  value;
    io_in_instrValid_15=value;
  endfunction

  function void get_io_in_pds_0_isRVCxxPfBDHPCKVf7;
    output logic  value;
    value=io_in_pds_0_isRVC;
  endfunction

  function void set_io_in_pds_0_isRVCxxPfBDHPCKVf7;
    input logic  value;
    io_in_pds_0_isRVC=value;
  endfunction

  function void get_io_in_pds_0_brTypexxPfBDHPCKVf7;
    output logic [1:0] value;
    value=io_in_pds_0_brType;
  endfunction

  function void set_io_in_pds_0_brTypexxPfBDHPCKVf7;
    input logic [1:0] value;
    io_in_pds_0_brType=value;
  endfunction

  function void get_io_in_pds_0_isRetxxPfBDHPCKVf7;
    output logic  value;
    value=io_in_pds_0_isRet;
  endfunction

  function void set_io_in_pds_0_isRetxxPfBDHPCKVf7;
    input logic  value;
    io_in_pds_0_isRet=value;
  endfunction

  function void get_io_in_pds_1_isRVCxxPfBDHPCKVf7;
    output logic  value;
    value=io_in_pds_1_isRVC;
  endfunction

  function void set_io_in_pds_1_isRVCxxPfBDHPCKVf7;
    input logic  value;
    io_in_pds_1_isRVC=value;
  endfunction

  function void get_io_in_pds_1_brTypexxPfBDHPCKVf7;
    output logic [1:0] value;
    value=io_in_pds_1_brType;
  endfunction

  function void set_io_in_pds_1_brTypexxPfBDHPCKVf7;
    input logic [1:0] value;
    io_in_pds_1_brType=value;
  endfunction

  function void get_io_in_pds_1_isRetxxPfBDHPCKVf7;
    output logic  value;
    value=io_in_pds_1_isRet;
  endfunction

  function void set_io_in_pds_1_isRetxxPfBDHPCKVf7;
    input logic  value;
    io_in_pds_1_isRet=value;
  endfunction

  function void get_io_in_pds_2_isRVCxxPfBDHPCKVf7;
    output logic  value;
    value=io_in_pds_2_isRVC;
  endfunction

  function void set_io_in_pds_2_isRVCxxPfBDHPCKVf7;
    input logic  value;
    io_in_pds_2_isRVC=value;
  endfunction

  function void get_io_in_pds_2_brTypexxPfBDHPCKVf7;
    output logic [1:0] value;
    value=io_in_pds_2_brType;
  endfunction

  function void set_io_in_pds_2_brTypexxPfBDHPCKVf7;
    input logic [1:0] value;
    io_in_pds_2_brType=value;
  endfunction

  function void get_io_in_pds_2_isRetxxPfBDHPCKVf7;
    output logic  value;
    value=io_in_pds_2_isRet;
  endfunction

  function void set_io_in_pds_2_isRetxxPfBDHPCKVf7;
    input logic  value;
    io_in_pds_2_isRet=value;
  endfunction

  function void get_io_in_pds_3_isRVCxxPfBDHPCKVf7;
    output logic  value;
    value=io_in_pds_3_isRVC;
  endfunction

  function void set_io_in_pds_3_isRVCxxPfBDHPCKVf7;
    input logic  value;
    io_in_pds_3_isRVC=value;
  endfunction

  function void get_io_in_pds_3_brTypexxPfBDHPCKVf7;
    output logic [1:0] value;
    value=io_in_pds_3_brType;
  endfunction

  function void set_io_in_pds_3_brTypexxPfBDHPCKVf7;
    input logic [1:0] value;
    io_in_pds_3_brType=value;
  endfunction

  function void get_io_in_pds_3_isRetxxPfBDHPCKVf7;
    output logic  value;
    value=io_in_pds_3_isRet;
  endfunction

  function void set_io_in_pds_3_isRetxxPfBDHPCKVf7;
    input logic  value;
    io_in_pds_3_isRet=value;
  endfunction

  function void get_io_in_pds_4_isRVCxxPfBDHPCKVf7;
    output logic  value;
    value=io_in_pds_4_isRVC;
  endfunction

  function void set_io_in_pds_4_isRVCxxPfBDHPCKVf7;
    input logic  value;
    io_in_pds_4_isRVC=value;
  endfunction

  function void get_io_in_pds_4_brTypexxPfBDHPCKVf7;
    output logic [1:0] value;
    value=io_in_pds_4_brType;
  endfunction

  function void set_io_in_pds_4_brTypexxPfBDHPCKVf7;
    input logic [1:0] value;
    io_in_pds_4_brType=value;
  endfunction

  function void get_io_in_pds_4_isRetxxPfBDHPCKVf7;
    output logic  value;
    value=io_in_pds_4_isRet;
  endfunction

  function void set_io_in_pds_4_isRetxxPfBDHPCKVf7;
    input logic  value;
    io_in_pds_4_isRet=value;
  endfunction

  function void get_io_in_pds_5_isRVCxxPfBDHPCKVf7;
    output logic  value;
    value=io_in_pds_5_isRVC;
  endfunction

  function void set_io_in_pds_5_isRVCxxPfBDHPCKVf7;
    input logic  value;
    io_in_pds_5_isRVC=value;
  endfunction

  function void get_io_in_pds_5_brTypexxPfBDHPCKVf7;
    output logic [1:0] value;
    value=io_in_pds_5_brType;
  endfunction

  function void set_io_in_pds_5_brTypexxPfBDHPCKVf7;
    input logic [1:0] value;
    io_in_pds_5_brType=value;
  endfunction

  function void get_io_in_pds_5_isRetxxPfBDHPCKVf7;
    output logic  value;
    value=io_in_pds_5_isRet;
  endfunction

  function void set_io_in_pds_5_isRetxxPfBDHPCKVf7;
    input logic  value;
    io_in_pds_5_isRet=value;
  endfunction

  function void get_io_in_pds_6_isRVCxxPfBDHPCKVf7;
    output logic  value;
    value=io_in_pds_6_isRVC;
  endfunction

  function void set_io_in_pds_6_isRVCxxPfBDHPCKVf7;
    input logic  value;
    io_in_pds_6_isRVC=value;
  endfunction

  function void get_io_in_pds_6_brTypexxPfBDHPCKVf7;
    output logic [1:0] value;
    value=io_in_pds_6_brType;
  endfunction

  function void set_io_in_pds_6_brTypexxPfBDHPCKVf7;
    input logic [1:0] value;
    io_in_pds_6_brType=value;
  endfunction

  function void get_io_in_pds_6_isRetxxPfBDHPCKVf7;
    output logic  value;
    value=io_in_pds_6_isRet;
  endfunction

  function void set_io_in_pds_6_isRetxxPfBDHPCKVf7;
    input logic  value;
    io_in_pds_6_isRet=value;
  endfunction

  function void get_io_in_pds_7_isRVCxxPfBDHPCKVf7;
    output logic  value;
    value=io_in_pds_7_isRVC;
  endfunction

  function void set_io_in_pds_7_isRVCxxPfBDHPCKVf7;
    input logic  value;
    io_in_pds_7_isRVC=value;
  endfunction

  function void get_io_in_pds_7_brTypexxPfBDHPCKVf7;
    output logic [1:0] value;
    value=io_in_pds_7_brType;
  endfunction

  function void set_io_in_pds_7_brTypexxPfBDHPCKVf7;
    input logic [1:0] value;
    io_in_pds_7_brType=value;
  endfunction

  function void get_io_in_pds_7_isRetxxPfBDHPCKVf7;
    output logic  value;
    value=io_in_pds_7_isRet;
  endfunction

  function void set_io_in_pds_7_isRetxxPfBDHPCKVf7;
    input logic  value;
    io_in_pds_7_isRet=value;
  endfunction

  function void get_io_in_pds_8_isRVCxxPfBDHPCKVf7;
    output logic  value;
    value=io_in_pds_8_isRVC;
  endfunction

  function void set_io_in_pds_8_isRVCxxPfBDHPCKVf7;
    input logic  value;
    io_in_pds_8_isRVC=value;
  endfunction

  function void get_io_in_pds_8_brTypexxPfBDHPCKVf7;
    output logic [1:0] value;
    value=io_in_pds_8_brType;
  endfunction

  function void set_io_in_pds_8_brTypexxPfBDHPCKVf7;
    input logic [1:0] value;
    io_in_pds_8_brType=value;
  endfunction

  function void get_io_in_pds_8_isRetxxPfBDHPCKVf7;
    output logic  value;
    value=io_in_pds_8_isRet;
  endfunction

  function void set_io_in_pds_8_isRetxxPfBDHPCKVf7;
    input logic  value;
    io_in_pds_8_isRet=value;
  endfunction

  function void get_io_in_pds_9_isRVCxxPfBDHPCKVf7;
    output logic  value;
    value=io_in_pds_9_isRVC;
  endfunction

  function void set_io_in_pds_9_isRVCxxPfBDHPCKVf7;
    input logic  value;
    io_in_pds_9_isRVC=value;
  endfunction

  function void get_io_in_pds_9_brTypexxPfBDHPCKVf7;
    output logic [1:0] value;
    value=io_in_pds_9_brType;
  endfunction

  function void set_io_in_pds_9_brTypexxPfBDHPCKVf7;
    input logic [1:0] value;
    io_in_pds_9_brType=value;
  endfunction

  function void get_io_in_pds_9_isRetxxPfBDHPCKVf7;
    output logic  value;
    value=io_in_pds_9_isRet;
  endfunction

  function void set_io_in_pds_9_isRetxxPfBDHPCKVf7;
    input logic  value;
    io_in_pds_9_isRet=value;
  endfunction

  function void get_io_in_pds_10_isRVCxxPfBDHPCKVf7;
    output logic  value;
    value=io_in_pds_10_isRVC;
  endfunction

  function void set_io_in_pds_10_isRVCxxPfBDHPCKVf7;
    input logic  value;
    io_in_pds_10_isRVC=value;
  endfunction

  function void get_io_in_pds_10_brTypexxPfBDHPCKVf7;
    output logic [1:0] value;
    value=io_in_pds_10_brType;
  endfunction

  function void set_io_in_pds_10_brTypexxPfBDHPCKVf7;
    input logic [1:0] value;
    io_in_pds_10_brType=value;
  endfunction

  function void get_io_in_pds_10_isRetxxPfBDHPCKVf7;
    output logic  value;
    value=io_in_pds_10_isRet;
  endfunction

  function void set_io_in_pds_10_isRetxxPfBDHPCKVf7;
    input logic  value;
    io_in_pds_10_isRet=value;
  endfunction

  function void get_io_in_pds_11_isRVCxxPfBDHPCKVf7;
    output logic  value;
    value=io_in_pds_11_isRVC;
  endfunction

  function void set_io_in_pds_11_isRVCxxPfBDHPCKVf7;
    input logic  value;
    io_in_pds_11_isRVC=value;
  endfunction

  function void get_io_in_pds_11_brTypexxPfBDHPCKVf7;
    output logic [1:0] value;
    value=io_in_pds_11_brType;
  endfunction

  function void set_io_in_pds_11_brTypexxPfBDHPCKVf7;
    input logic [1:0] value;
    io_in_pds_11_brType=value;
  endfunction

  function void get_io_in_pds_11_isRetxxPfBDHPCKVf7;
    output logic  value;
    value=io_in_pds_11_isRet;
  endfunction

  function void set_io_in_pds_11_isRetxxPfBDHPCKVf7;
    input logic  value;
    io_in_pds_11_isRet=value;
  endfunction

  function void get_io_in_pds_12_isRVCxxPfBDHPCKVf7;
    output logic  value;
    value=io_in_pds_12_isRVC;
  endfunction

  function void set_io_in_pds_12_isRVCxxPfBDHPCKVf7;
    input logic  value;
    io_in_pds_12_isRVC=value;
  endfunction

  function void get_io_in_pds_12_brTypexxPfBDHPCKVf7;
    output logic [1:0] value;
    value=io_in_pds_12_brType;
  endfunction

  function void set_io_in_pds_12_brTypexxPfBDHPCKVf7;
    input logic [1:0] value;
    io_in_pds_12_brType=value;
  endfunction

  function void get_io_in_pds_12_isRetxxPfBDHPCKVf7;
    output logic  value;
    value=io_in_pds_12_isRet;
  endfunction

  function void set_io_in_pds_12_isRetxxPfBDHPCKVf7;
    input logic  value;
    io_in_pds_12_isRet=value;
  endfunction

  function void get_io_in_pds_13_isRVCxxPfBDHPCKVf7;
    output logic  value;
    value=io_in_pds_13_isRVC;
  endfunction

  function void set_io_in_pds_13_isRVCxxPfBDHPCKVf7;
    input logic  value;
    io_in_pds_13_isRVC=value;
  endfunction

  function void get_io_in_pds_13_brTypexxPfBDHPCKVf7;
    output logic [1:0] value;
    value=io_in_pds_13_brType;
  endfunction

  function void set_io_in_pds_13_brTypexxPfBDHPCKVf7;
    input logic [1:0] value;
    io_in_pds_13_brType=value;
  endfunction

  function void get_io_in_pds_13_isRetxxPfBDHPCKVf7;
    output logic  value;
    value=io_in_pds_13_isRet;
  endfunction

  function void set_io_in_pds_13_isRetxxPfBDHPCKVf7;
    input logic  value;
    io_in_pds_13_isRet=value;
  endfunction

  function void get_io_in_pds_14_isRVCxxPfBDHPCKVf7;
    output logic  value;
    value=io_in_pds_14_isRVC;
  endfunction

  function void set_io_in_pds_14_isRVCxxPfBDHPCKVf7;
    input logic  value;
    io_in_pds_14_isRVC=value;
  endfunction

  function void get_io_in_pds_14_brTypexxPfBDHPCKVf7;
    output logic [1:0] value;
    value=io_in_pds_14_brType;
  endfunction

  function void set_io_in_pds_14_brTypexxPfBDHPCKVf7;
    input logic [1:0] value;
    io_in_pds_14_brType=value;
  endfunction

  function void get_io_in_pds_14_isRetxxPfBDHPCKVf7;
    output logic  value;
    value=io_in_pds_14_isRet;
  endfunction

  function void set_io_in_pds_14_isRetxxPfBDHPCKVf7;
    input logic  value;
    io_in_pds_14_isRet=value;
  endfunction

  function void get_io_in_pds_15_isRVCxxPfBDHPCKVf7;
    output logic  value;
    value=io_in_pds_15_isRVC;
  endfunction

  function void set_io_in_pds_15_isRVCxxPfBDHPCKVf7;
    input logic  value;
    io_in_pds_15_isRVC=value;
  endfunction

  function void get_io_in_pds_15_brTypexxPfBDHPCKVf7;
    output logic [1:0] value;
    value=io_in_pds_15_brType;
  endfunction

  function void set_io_in_pds_15_brTypexxPfBDHPCKVf7;
    input logic [1:0] value;
    io_in_pds_15_brType=value;
  endfunction

  function void get_io_in_pds_15_isRetxxPfBDHPCKVf7;
    output logic  value;
    value=io_in_pds_15_isRet;
  endfunction

  function void set_io_in_pds_15_isRetxxPfBDHPCKVf7;
    input logic  value;
    io_in_pds_15_isRet=value;
  endfunction

  function void get_io_in_pc_0xxPfBDHPCKVf7;
    output logic [49:0] value;
    value=io_in_pc_0;
  endfunction

  function void set_io_in_pc_0xxPfBDHPCKVf7;
    input logic [49:0] value;
    io_in_pc_0=value;
  endfunction

  function void get_io_in_pc_1xxPfBDHPCKVf7;
    output logic [49:0] value;
    value=io_in_pc_1;
  endfunction

  function void set_io_in_pc_1xxPfBDHPCKVf7;
    input logic [49:0] value;
    io_in_pc_1=value;
  endfunction

  function void get_io_in_pc_2xxPfBDHPCKVf7;
    output logic [49:0] value;
    value=io_in_pc_2;
  endfunction

  function void set_io_in_pc_2xxPfBDHPCKVf7;
    input logic [49:0] value;
    io_in_pc_2=value;
  endfunction

  function void get_io_in_pc_3xxPfBDHPCKVf7;
    output logic [49:0] value;
    value=io_in_pc_3;
  endfunction

  function void set_io_in_pc_3xxPfBDHPCKVf7;
    input logic [49:0] value;
    io_in_pc_3=value;
  endfunction

  function void get_io_in_pc_4xxPfBDHPCKVf7;
    output logic [49:0] value;
    value=io_in_pc_4;
  endfunction

  function void set_io_in_pc_4xxPfBDHPCKVf7;
    input logic [49:0] value;
    io_in_pc_4=value;
  endfunction

  function void get_io_in_pc_5xxPfBDHPCKVf7;
    output logic [49:0] value;
    value=io_in_pc_5;
  endfunction

  function void set_io_in_pc_5xxPfBDHPCKVf7;
    input logic [49:0] value;
    io_in_pc_5=value;
  endfunction

  function void get_io_in_pc_6xxPfBDHPCKVf7;
    output logic [49:0] value;
    value=io_in_pc_6;
  endfunction

  function void set_io_in_pc_6xxPfBDHPCKVf7;
    input logic [49:0] value;
    io_in_pc_6=value;
  endfunction

  function void get_io_in_pc_7xxPfBDHPCKVf7;
    output logic [49:0] value;
    value=io_in_pc_7;
  endfunction

  function void set_io_in_pc_7xxPfBDHPCKVf7;
    input logic [49:0] value;
    io_in_pc_7=value;
  endfunction

  function void get_io_in_pc_8xxPfBDHPCKVf7;
    output logic [49:0] value;
    value=io_in_pc_8;
  endfunction

  function void set_io_in_pc_8xxPfBDHPCKVf7;
    input logic [49:0] value;
    io_in_pc_8=value;
  endfunction

  function void get_io_in_pc_9xxPfBDHPCKVf7;
    output logic [49:0] value;
    value=io_in_pc_9;
  endfunction

  function void set_io_in_pc_9xxPfBDHPCKVf7;
    input logic [49:0] value;
    io_in_pc_9=value;
  endfunction

  function void get_io_in_pc_10xxPfBDHPCKVf7;
    output logic [49:0] value;
    value=io_in_pc_10;
  endfunction

  function void set_io_in_pc_10xxPfBDHPCKVf7;
    input logic [49:0] value;
    io_in_pc_10=value;
  endfunction

  function void get_io_in_pc_11xxPfBDHPCKVf7;
    output logic [49:0] value;
    value=io_in_pc_11;
  endfunction

  function void set_io_in_pc_11xxPfBDHPCKVf7;
    input logic [49:0] value;
    io_in_pc_11=value;
  endfunction

  function void get_io_in_pc_12xxPfBDHPCKVf7;
    output logic [49:0] value;
    value=io_in_pc_12;
  endfunction

  function void set_io_in_pc_12xxPfBDHPCKVf7;
    input logic [49:0] value;
    io_in_pc_12=value;
  endfunction

  function void get_io_in_pc_13xxPfBDHPCKVf7;
    output logic [49:0] value;
    value=io_in_pc_13;
  endfunction

  function void set_io_in_pc_13xxPfBDHPCKVf7;
    input logic [49:0] value;
    io_in_pc_13=value;
  endfunction

  function void get_io_in_pc_14xxPfBDHPCKVf7;
    output logic [49:0] value;
    value=io_in_pc_14;
  endfunction

  function void set_io_in_pc_14xxPfBDHPCKVf7;
    input logic [49:0] value;
    io_in_pc_14=value;
  endfunction

  function void get_io_in_pc_15xxPfBDHPCKVf7;
    output logic [49:0] value;
    value=io_in_pc_15;
  endfunction

  function void set_io_in_pc_15xxPfBDHPCKVf7;
    input logic [49:0] value;
    io_in_pc_15=value;
  endfunction

  function void get_io_in_fire_inxxPfBDHPCKVf7;
    output logic  value;
    value=io_in_fire_in;
  endfunction

  function void set_io_in_fire_inxxPfBDHPCKVf7;
    input logic  value;
    io_in_fire_in=value;
  endfunction

  function void get_io_out_stage1Out_fixedRange_0xxPfBDHPCKVf7;
    output logic  value;
    value=io_out_stage1Out_fixedRange_0;
  endfunction

  function void set_io_out_stage1Out_fixedRange_0xxPfBDHPCKVf7;
    input logic  value;
    io_out_stage1Out_fixedRange_0=value;
  endfunction

  function void get_io_out_stage1Out_fixedRange_1xxPfBDHPCKVf7;
    output logic  value;
    value=io_out_stage1Out_fixedRange_1;
  endfunction

  function void set_io_out_stage1Out_fixedRange_1xxPfBDHPCKVf7;
    input logic  value;
    io_out_stage1Out_fixedRange_1=value;
  endfunction

  function void get_io_out_stage1Out_fixedRange_2xxPfBDHPCKVf7;
    output logic  value;
    value=io_out_stage1Out_fixedRange_2;
  endfunction

  function void set_io_out_stage1Out_fixedRange_2xxPfBDHPCKVf7;
    input logic  value;
    io_out_stage1Out_fixedRange_2=value;
  endfunction

  function void get_io_out_stage1Out_fixedRange_3xxPfBDHPCKVf7;
    output logic  value;
    value=io_out_stage1Out_fixedRange_3;
  endfunction

  function void set_io_out_stage1Out_fixedRange_3xxPfBDHPCKVf7;
    input logic  value;
    io_out_stage1Out_fixedRange_3=value;
  endfunction

  function void get_io_out_stage1Out_fixedRange_4xxPfBDHPCKVf7;
    output logic  value;
    value=io_out_stage1Out_fixedRange_4;
  endfunction

  function void set_io_out_stage1Out_fixedRange_4xxPfBDHPCKVf7;
    input logic  value;
    io_out_stage1Out_fixedRange_4=value;
  endfunction

  function void get_io_out_stage1Out_fixedRange_5xxPfBDHPCKVf7;
    output logic  value;
    value=io_out_stage1Out_fixedRange_5;
  endfunction

  function void set_io_out_stage1Out_fixedRange_5xxPfBDHPCKVf7;
    input logic  value;
    io_out_stage1Out_fixedRange_5=value;
  endfunction

  function void get_io_out_stage1Out_fixedRange_6xxPfBDHPCKVf7;
    output logic  value;
    value=io_out_stage1Out_fixedRange_6;
  endfunction

  function void set_io_out_stage1Out_fixedRange_6xxPfBDHPCKVf7;
    input logic  value;
    io_out_stage1Out_fixedRange_6=value;
  endfunction

  function void get_io_out_stage1Out_fixedRange_7xxPfBDHPCKVf7;
    output logic  value;
    value=io_out_stage1Out_fixedRange_7;
  endfunction

  function void set_io_out_stage1Out_fixedRange_7xxPfBDHPCKVf7;
    input logic  value;
    io_out_stage1Out_fixedRange_7=value;
  endfunction

  function void get_io_out_stage1Out_fixedRange_8xxPfBDHPCKVf7;
    output logic  value;
    value=io_out_stage1Out_fixedRange_8;
  endfunction

  function void set_io_out_stage1Out_fixedRange_8xxPfBDHPCKVf7;
    input logic  value;
    io_out_stage1Out_fixedRange_8=value;
  endfunction

  function void get_io_out_stage1Out_fixedRange_9xxPfBDHPCKVf7;
    output logic  value;
    value=io_out_stage1Out_fixedRange_9;
  endfunction

  function void set_io_out_stage1Out_fixedRange_9xxPfBDHPCKVf7;
    input logic  value;
    io_out_stage1Out_fixedRange_9=value;
  endfunction

  function void get_io_out_stage1Out_fixedRange_10xxPfBDHPCKVf7;
    output logic  value;
    value=io_out_stage1Out_fixedRange_10;
  endfunction

  function void set_io_out_stage1Out_fixedRange_10xxPfBDHPCKVf7;
    input logic  value;
    io_out_stage1Out_fixedRange_10=value;
  endfunction

  function void get_io_out_stage1Out_fixedRange_11xxPfBDHPCKVf7;
    output logic  value;
    value=io_out_stage1Out_fixedRange_11;
  endfunction

  function void set_io_out_stage1Out_fixedRange_11xxPfBDHPCKVf7;
    input logic  value;
    io_out_stage1Out_fixedRange_11=value;
  endfunction

  function void get_io_out_stage1Out_fixedRange_12xxPfBDHPCKVf7;
    output logic  value;
    value=io_out_stage1Out_fixedRange_12;
  endfunction

  function void set_io_out_stage1Out_fixedRange_12xxPfBDHPCKVf7;
    input logic  value;
    io_out_stage1Out_fixedRange_12=value;
  endfunction

  function void get_io_out_stage1Out_fixedRange_13xxPfBDHPCKVf7;
    output logic  value;
    value=io_out_stage1Out_fixedRange_13;
  endfunction

  function void set_io_out_stage1Out_fixedRange_13xxPfBDHPCKVf7;
    input logic  value;
    io_out_stage1Out_fixedRange_13=value;
  endfunction

  function void get_io_out_stage1Out_fixedRange_14xxPfBDHPCKVf7;
    output logic  value;
    value=io_out_stage1Out_fixedRange_14;
  endfunction

  function void set_io_out_stage1Out_fixedRange_14xxPfBDHPCKVf7;
    input logic  value;
    io_out_stage1Out_fixedRange_14=value;
  endfunction

  function void get_io_out_stage1Out_fixedRange_15xxPfBDHPCKVf7;
    output logic  value;
    value=io_out_stage1Out_fixedRange_15;
  endfunction

  function void set_io_out_stage1Out_fixedRange_15xxPfBDHPCKVf7;
    input logic  value;
    io_out_stage1Out_fixedRange_15=value;
  endfunction

  function void get_io_out_stage1Out_fixedTaken_0xxPfBDHPCKVf7;
    output logic  value;
    value=io_out_stage1Out_fixedTaken_0;
  endfunction

  function void set_io_out_stage1Out_fixedTaken_0xxPfBDHPCKVf7;
    input logic  value;
    io_out_stage1Out_fixedTaken_0=value;
  endfunction

  function void get_io_out_stage1Out_fixedTaken_1xxPfBDHPCKVf7;
    output logic  value;
    value=io_out_stage1Out_fixedTaken_1;
  endfunction

  function void set_io_out_stage1Out_fixedTaken_1xxPfBDHPCKVf7;
    input logic  value;
    io_out_stage1Out_fixedTaken_1=value;
  endfunction

  function void get_io_out_stage1Out_fixedTaken_2xxPfBDHPCKVf7;
    output logic  value;
    value=io_out_stage1Out_fixedTaken_2;
  endfunction

  function void set_io_out_stage1Out_fixedTaken_2xxPfBDHPCKVf7;
    input logic  value;
    io_out_stage1Out_fixedTaken_2=value;
  endfunction

  function void get_io_out_stage1Out_fixedTaken_3xxPfBDHPCKVf7;
    output logic  value;
    value=io_out_stage1Out_fixedTaken_3;
  endfunction

  function void set_io_out_stage1Out_fixedTaken_3xxPfBDHPCKVf7;
    input logic  value;
    io_out_stage1Out_fixedTaken_3=value;
  endfunction

  function void get_io_out_stage1Out_fixedTaken_4xxPfBDHPCKVf7;
    output logic  value;
    value=io_out_stage1Out_fixedTaken_4;
  endfunction

  function void set_io_out_stage1Out_fixedTaken_4xxPfBDHPCKVf7;
    input logic  value;
    io_out_stage1Out_fixedTaken_4=value;
  endfunction

  function void get_io_out_stage1Out_fixedTaken_5xxPfBDHPCKVf7;
    output logic  value;
    value=io_out_stage1Out_fixedTaken_5;
  endfunction

  function void set_io_out_stage1Out_fixedTaken_5xxPfBDHPCKVf7;
    input logic  value;
    io_out_stage1Out_fixedTaken_5=value;
  endfunction

  function void get_io_out_stage1Out_fixedTaken_6xxPfBDHPCKVf7;
    output logic  value;
    value=io_out_stage1Out_fixedTaken_6;
  endfunction

  function void set_io_out_stage1Out_fixedTaken_6xxPfBDHPCKVf7;
    input logic  value;
    io_out_stage1Out_fixedTaken_6=value;
  endfunction

  function void get_io_out_stage1Out_fixedTaken_7xxPfBDHPCKVf7;
    output logic  value;
    value=io_out_stage1Out_fixedTaken_7;
  endfunction

  function void set_io_out_stage1Out_fixedTaken_7xxPfBDHPCKVf7;
    input logic  value;
    io_out_stage1Out_fixedTaken_7=value;
  endfunction

  function void get_io_out_stage1Out_fixedTaken_8xxPfBDHPCKVf7;
    output logic  value;
    value=io_out_stage1Out_fixedTaken_8;
  endfunction

  function void set_io_out_stage1Out_fixedTaken_8xxPfBDHPCKVf7;
    input logic  value;
    io_out_stage1Out_fixedTaken_8=value;
  endfunction

  function void get_io_out_stage1Out_fixedTaken_9xxPfBDHPCKVf7;
    output logic  value;
    value=io_out_stage1Out_fixedTaken_9;
  endfunction

  function void set_io_out_stage1Out_fixedTaken_9xxPfBDHPCKVf7;
    input logic  value;
    io_out_stage1Out_fixedTaken_9=value;
  endfunction

  function void get_io_out_stage1Out_fixedTaken_10xxPfBDHPCKVf7;
    output logic  value;
    value=io_out_stage1Out_fixedTaken_10;
  endfunction

  function void set_io_out_stage1Out_fixedTaken_10xxPfBDHPCKVf7;
    input logic  value;
    io_out_stage1Out_fixedTaken_10=value;
  endfunction

  function void get_io_out_stage1Out_fixedTaken_11xxPfBDHPCKVf7;
    output logic  value;
    value=io_out_stage1Out_fixedTaken_11;
  endfunction

  function void set_io_out_stage1Out_fixedTaken_11xxPfBDHPCKVf7;
    input logic  value;
    io_out_stage1Out_fixedTaken_11=value;
  endfunction

  function void get_io_out_stage1Out_fixedTaken_12xxPfBDHPCKVf7;
    output logic  value;
    value=io_out_stage1Out_fixedTaken_12;
  endfunction

  function void set_io_out_stage1Out_fixedTaken_12xxPfBDHPCKVf7;
    input logic  value;
    io_out_stage1Out_fixedTaken_12=value;
  endfunction

  function void get_io_out_stage1Out_fixedTaken_13xxPfBDHPCKVf7;
    output logic  value;
    value=io_out_stage1Out_fixedTaken_13;
  endfunction

  function void set_io_out_stage1Out_fixedTaken_13xxPfBDHPCKVf7;
    input logic  value;
    io_out_stage1Out_fixedTaken_13=value;
  endfunction

  function void get_io_out_stage1Out_fixedTaken_14xxPfBDHPCKVf7;
    output logic  value;
    value=io_out_stage1Out_fixedTaken_14;
  endfunction

  function void set_io_out_stage1Out_fixedTaken_14xxPfBDHPCKVf7;
    input logic  value;
    io_out_stage1Out_fixedTaken_14=value;
  endfunction

  function void get_io_out_stage1Out_fixedTaken_15xxPfBDHPCKVf7;
    output logic  value;
    value=io_out_stage1Out_fixedTaken_15;
  endfunction

  function void set_io_out_stage1Out_fixedTaken_15xxPfBDHPCKVf7;
    input logic  value;
    io_out_stage1Out_fixedTaken_15=value;
  endfunction

  function void get_io_out_stage2Out_fixedTarget_0xxPfBDHPCKVf7;
    output logic [49:0] value;
    value=io_out_stage2Out_fixedTarget_0;
  endfunction

  function void set_io_out_stage2Out_fixedTarget_0xxPfBDHPCKVf7;
    input logic [49:0] value;
    io_out_stage2Out_fixedTarget_0=value;
  endfunction

  function void get_io_out_stage2Out_fixedTarget_1xxPfBDHPCKVf7;
    output logic [49:0] value;
    value=io_out_stage2Out_fixedTarget_1;
  endfunction

  function void set_io_out_stage2Out_fixedTarget_1xxPfBDHPCKVf7;
    input logic [49:0] value;
    io_out_stage2Out_fixedTarget_1=value;
  endfunction

  function void get_io_out_stage2Out_fixedTarget_2xxPfBDHPCKVf7;
    output logic [49:0] value;
    value=io_out_stage2Out_fixedTarget_2;
  endfunction

  function void set_io_out_stage2Out_fixedTarget_2xxPfBDHPCKVf7;
    input logic [49:0] value;
    io_out_stage2Out_fixedTarget_2=value;
  endfunction

  function void get_io_out_stage2Out_fixedTarget_3xxPfBDHPCKVf7;
    output logic [49:0] value;
    value=io_out_stage2Out_fixedTarget_3;
  endfunction

  function void set_io_out_stage2Out_fixedTarget_3xxPfBDHPCKVf7;
    input logic [49:0] value;
    io_out_stage2Out_fixedTarget_3=value;
  endfunction

  function void get_io_out_stage2Out_fixedTarget_4xxPfBDHPCKVf7;
    output logic [49:0] value;
    value=io_out_stage2Out_fixedTarget_4;
  endfunction

  function void set_io_out_stage2Out_fixedTarget_4xxPfBDHPCKVf7;
    input logic [49:0] value;
    io_out_stage2Out_fixedTarget_4=value;
  endfunction

  function void get_io_out_stage2Out_fixedTarget_5xxPfBDHPCKVf7;
    output logic [49:0] value;
    value=io_out_stage2Out_fixedTarget_5;
  endfunction

  function void set_io_out_stage2Out_fixedTarget_5xxPfBDHPCKVf7;
    input logic [49:0] value;
    io_out_stage2Out_fixedTarget_5=value;
  endfunction

  function void get_io_out_stage2Out_fixedTarget_6xxPfBDHPCKVf7;
    output logic [49:0] value;
    value=io_out_stage2Out_fixedTarget_6;
  endfunction

  function void set_io_out_stage2Out_fixedTarget_6xxPfBDHPCKVf7;
    input logic [49:0] value;
    io_out_stage2Out_fixedTarget_6=value;
  endfunction

  function void get_io_out_stage2Out_fixedTarget_7xxPfBDHPCKVf7;
    output logic [49:0] value;
    value=io_out_stage2Out_fixedTarget_7;
  endfunction

  function void set_io_out_stage2Out_fixedTarget_7xxPfBDHPCKVf7;
    input logic [49:0] value;
    io_out_stage2Out_fixedTarget_7=value;
  endfunction

  function void get_io_out_stage2Out_fixedTarget_8xxPfBDHPCKVf7;
    output logic [49:0] value;
    value=io_out_stage2Out_fixedTarget_8;
  endfunction

  function void set_io_out_stage2Out_fixedTarget_8xxPfBDHPCKVf7;
    input logic [49:0] value;
    io_out_stage2Out_fixedTarget_8=value;
  endfunction

  function void get_io_out_stage2Out_fixedTarget_9xxPfBDHPCKVf7;
    output logic [49:0] value;
    value=io_out_stage2Out_fixedTarget_9;
  endfunction

  function void set_io_out_stage2Out_fixedTarget_9xxPfBDHPCKVf7;
    input logic [49:0] value;
    io_out_stage2Out_fixedTarget_9=value;
  endfunction

  function void get_io_out_stage2Out_fixedTarget_10xxPfBDHPCKVf7;
    output logic [49:0] value;
    value=io_out_stage2Out_fixedTarget_10;
  endfunction

  function void set_io_out_stage2Out_fixedTarget_10xxPfBDHPCKVf7;
    input logic [49:0] value;
    io_out_stage2Out_fixedTarget_10=value;
  endfunction

  function void get_io_out_stage2Out_fixedTarget_11xxPfBDHPCKVf7;
    output logic [49:0] value;
    value=io_out_stage2Out_fixedTarget_11;
  endfunction

  function void set_io_out_stage2Out_fixedTarget_11xxPfBDHPCKVf7;
    input logic [49:0] value;
    io_out_stage2Out_fixedTarget_11=value;
  endfunction

  function void get_io_out_stage2Out_fixedTarget_12xxPfBDHPCKVf7;
    output logic [49:0] value;
    value=io_out_stage2Out_fixedTarget_12;
  endfunction

  function void set_io_out_stage2Out_fixedTarget_12xxPfBDHPCKVf7;
    input logic [49:0] value;
    io_out_stage2Out_fixedTarget_12=value;
  endfunction

  function void get_io_out_stage2Out_fixedTarget_13xxPfBDHPCKVf7;
    output logic [49:0] value;
    value=io_out_stage2Out_fixedTarget_13;
  endfunction

  function void set_io_out_stage2Out_fixedTarget_13xxPfBDHPCKVf7;
    input logic [49:0] value;
    io_out_stage2Out_fixedTarget_13=value;
  endfunction

  function void get_io_out_stage2Out_fixedTarget_14xxPfBDHPCKVf7;
    output logic [49:0] value;
    value=io_out_stage2Out_fixedTarget_14;
  endfunction

  function void set_io_out_stage2Out_fixedTarget_14xxPfBDHPCKVf7;
    input logic [49:0] value;
    io_out_stage2Out_fixedTarget_14=value;
  endfunction

  function void get_io_out_stage2Out_fixedTarget_15xxPfBDHPCKVf7;
    output logic [49:0] value;
    value=io_out_stage2Out_fixedTarget_15;
  endfunction

  function void set_io_out_stage2Out_fixedTarget_15xxPfBDHPCKVf7;
    input logic [49:0] value;
    io_out_stage2Out_fixedTarget_15=value;
  endfunction

  function void get_io_out_stage2Out_jalTarget_0xxPfBDHPCKVf7;
    output logic [49:0] value;
    value=io_out_stage2Out_jalTarget_0;
  endfunction

  function void set_io_out_stage2Out_jalTarget_0xxPfBDHPCKVf7;
    input logic [49:0] value;
    io_out_stage2Out_jalTarget_0=value;
  endfunction

  function void get_io_out_stage2Out_jalTarget_1xxPfBDHPCKVf7;
    output logic [49:0] value;
    value=io_out_stage2Out_jalTarget_1;
  endfunction

  function void set_io_out_stage2Out_jalTarget_1xxPfBDHPCKVf7;
    input logic [49:0] value;
    io_out_stage2Out_jalTarget_1=value;
  endfunction

  function void get_io_out_stage2Out_jalTarget_2xxPfBDHPCKVf7;
    output logic [49:0] value;
    value=io_out_stage2Out_jalTarget_2;
  endfunction

  function void set_io_out_stage2Out_jalTarget_2xxPfBDHPCKVf7;
    input logic [49:0] value;
    io_out_stage2Out_jalTarget_2=value;
  endfunction

  function void get_io_out_stage2Out_jalTarget_3xxPfBDHPCKVf7;
    output logic [49:0] value;
    value=io_out_stage2Out_jalTarget_3;
  endfunction

  function void set_io_out_stage2Out_jalTarget_3xxPfBDHPCKVf7;
    input logic [49:0] value;
    io_out_stage2Out_jalTarget_3=value;
  endfunction

  function void get_io_out_stage2Out_jalTarget_4xxPfBDHPCKVf7;
    output logic [49:0] value;
    value=io_out_stage2Out_jalTarget_4;
  endfunction

  function void set_io_out_stage2Out_jalTarget_4xxPfBDHPCKVf7;
    input logic [49:0] value;
    io_out_stage2Out_jalTarget_4=value;
  endfunction

  function void get_io_out_stage2Out_jalTarget_5xxPfBDHPCKVf7;
    output logic [49:0] value;
    value=io_out_stage2Out_jalTarget_5;
  endfunction

  function void set_io_out_stage2Out_jalTarget_5xxPfBDHPCKVf7;
    input logic [49:0] value;
    io_out_stage2Out_jalTarget_5=value;
  endfunction

  function void get_io_out_stage2Out_jalTarget_6xxPfBDHPCKVf7;
    output logic [49:0] value;
    value=io_out_stage2Out_jalTarget_6;
  endfunction

  function void set_io_out_stage2Out_jalTarget_6xxPfBDHPCKVf7;
    input logic [49:0] value;
    io_out_stage2Out_jalTarget_6=value;
  endfunction

  function void get_io_out_stage2Out_jalTarget_7xxPfBDHPCKVf7;
    output logic [49:0] value;
    value=io_out_stage2Out_jalTarget_7;
  endfunction

  function void set_io_out_stage2Out_jalTarget_7xxPfBDHPCKVf7;
    input logic [49:0] value;
    io_out_stage2Out_jalTarget_7=value;
  endfunction

  function void get_io_out_stage2Out_jalTarget_8xxPfBDHPCKVf7;
    output logic [49:0] value;
    value=io_out_stage2Out_jalTarget_8;
  endfunction

  function void set_io_out_stage2Out_jalTarget_8xxPfBDHPCKVf7;
    input logic [49:0] value;
    io_out_stage2Out_jalTarget_8=value;
  endfunction

  function void get_io_out_stage2Out_jalTarget_9xxPfBDHPCKVf7;
    output logic [49:0] value;
    value=io_out_stage2Out_jalTarget_9;
  endfunction

  function void set_io_out_stage2Out_jalTarget_9xxPfBDHPCKVf7;
    input logic [49:0] value;
    io_out_stage2Out_jalTarget_9=value;
  endfunction

  function void get_io_out_stage2Out_jalTarget_10xxPfBDHPCKVf7;
    output logic [49:0] value;
    value=io_out_stage2Out_jalTarget_10;
  endfunction

  function void set_io_out_stage2Out_jalTarget_10xxPfBDHPCKVf7;
    input logic [49:0] value;
    io_out_stage2Out_jalTarget_10=value;
  endfunction

  function void get_io_out_stage2Out_jalTarget_11xxPfBDHPCKVf7;
    output logic [49:0] value;
    value=io_out_stage2Out_jalTarget_11;
  endfunction

  function void set_io_out_stage2Out_jalTarget_11xxPfBDHPCKVf7;
    input logic [49:0] value;
    io_out_stage2Out_jalTarget_11=value;
  endfunction

  function void get_io_out_stage2Out_jalTarget_12xxPfBDHPCKVf7;
    output logic [49:0] value;
    value=io_out_stage2Out_jalTarget_12;
  endfunction

  function void set_io_out_stage2Out_jalTarget_12xxPfBDHPCKVf7;
    input logic [49:0] value;
    io_out_stage2Out_jalTarget_12=value;
  endfunction

  function void get_io_out_stage2Out_jalTarget_13xxPfBDHPCKVf7;
    output logic [49:0] value;
    value=io_out_stage2Out_jalTarget_13;
  endfunction

  function void set_io_out_stage2Out_jalTarget_13xxPfBDHPCKVf7;
    input logic [49:0] value;
    io_out_stage2Out_jalTarget_13=value;
  endfunction

  function void get_io_out_stage2Out_jalTarget_14xxPfBDHPCKVf7;
    output logic [49:0] value;
    value=io_out_stage2Out_jalTarget_14;
  endfunction

  function void set_io_out_stage2Out_jalTarget_14xxPfBDHPCKVf7;
    input logic [49:0] value;
    io_out_stage2Out_jalTarget_14=value;
  endfunction

  function void get_io_out_stage2Out_jalTarget_15xxPfBDHPCKVf7;
    output logic [49:0] value;
    value=io_out_stage2Out_jalTarget_15;
  endfunction

  function void set_io_out_stage2Out_jalTarget_15xxPfBDHPCKVf7;
    input logic [49:0] value;
    io_out_stage2Out_jalTarget_15=value;
  endfunction

  function void get_io_out_stage2Out_fixedMissPred_0xxPfBDHPCKVf7;
    output logic  value;
    value=io_out_stage2Out_fixedMissPred_0;
  endfunction

  function void set_io_out_stage2Out_fixedMissPred_0xxPfBDHPCKVf7;
    input logic  value;
    io_out_stage2Out_fixedMissPred_0=value;
  endfunction

  function void get_io_out_stage2Out_fixedMissPred_1xxPfBDHPCKVf7;
    output logic  value;
    value=io_out_stage2Out_fixedMissPred_1;
  endfunction

  function void set_io_out_stage2Out_fixedMissPred_1xxPfBDHPCKVf7;
    input logic  value;
    io_out_stage2Out_fixedMissPred_1=value;
  endfunction

  function void get_io_out_stage2Out_fixedMissPred_2xxPfBDHPCKVf7;
    output logic  value;
    value=io_out_stage2Out_fixedMissPred_2;
  endfunction

  function void set_io_out_stage2Out_fixedMissPred_2xxPfBDHPCKVf7;
    input logic  value;
    io_out_stage2Out_fixedMissPred_2=value;
  endfunction

  function void get_io_out_stage2Out_fixedMissPred_3xxPfBDHPCKVf7;
    output logic  value;
    value=io_out_stage2Out_fixedMissPred_3;
  endfunction

  function void set_io_out_stage2Out_fixedMissPred_3xxPfBDHPCKVf7;
    input logic  value;
    io_out_stage2Out_fixedMissPred_3=value;
  endfunction

  function void get_io_out_stage2Out_fixedMissPred_4xxPfBDHPCKVf7;
    output logic  value;
    value=io_out_stage2Out_fixedMissPred_4;
  endfunction

  function void set_io_out_stage2Out_fixedMissPred_4xxPfBDHPCKVf7;
    input logic  value;
    io_out_stage2Out_fixedMissPred_4=value;
  endfunction

  function void get_io_out_stage2Out_fixedMissPred_5xxPfBDHPCKVf7;
    output logic  value;
    value=io_out_stage2Out_fixedMissPred_5;
  endfunction

  function void set_io_out_stage2Out_fixedMissPred_5xxPfBDHPCKVf7;
    input logic  value;
    io_out_stage2Out_fixedMissPred_5=value;
  endfunction

  function void get_io_out_stage2Out_fixedMissPred_6xxPfBDHPCKVf7;
    output logic  value;
    value=io_out_stage2Out_fixedMissPred_6;
  endfunction

  function void set_io_out_stage2Out_fixedMissPred_6xxPfBDHPCKVf7;
    input logic  value;
    io_out_stage2Out_fixedMissPred_6=value;
  endfunction

  function void get_io_out_stage2Out_fixedMissPred_7xxPfBDHPCKVf7;
    output logic  value;
    value=io_out_stage2Out_fixedMissPred_7;
  endfunction

  function void set_io_out_stage2Out_fixedMissPred_7xxPfBDHPCKVf7;
    input logic  value;
    io_out_stage2Out_fixedMissPred_7=value;
  endfunction

  function void get_io_out_stage2Out_fixedMissPred_8xxPfBDHPCKVf7;
    output logic  value;
    value=io_out_stage2Out_fixedMissPred_8;
  endfunction

  function void set_io_out_stage2Out_fixedMissPred_8xxPfBDHPCKVf7;
    input logic  value;
    io_out_stage2Out_fixedMissPred_8=value;
  endfunction

  function void get_io_out_stage2Out_fixedMissPred_9xxPfBDHPCKVf7;
    output logic  value;
    value=io_out_stage2Out_fixedMissPred_9;
  endfunction

  function void set_io_out_stage2Out_fixedMissPred_9xxPfBDHPCKVf7;
    input logic  value;
    io_out_stage2Out_fixedMissPred_9=value;
  endfunction

  function void get_io_out_stage2Out_fixedMissPred_10xxPfBDHPCKVf7;
    output logic  value;
    value=io_out_stage2Out_fixedMissPred_10;
  endfunction

  function void set_io_out_stage2Out_fixedMissPred_10xxPfBDHPCKVf7;
    input logic  value;
    io_out_stage2Out_fixedMissPred_10=value;
  endfunction

  function void get_io_out_stage2Out_fixedMissPred_11xxPfBDHPCKVf7;
    output logic  value;
    value=io_out_stage2Out_fixedMissPred_11;
  endfunction

  function void set_io_out_stage2Out_fixedMissPred_11xxPfBDHPCKVf7;
    input logic  value;
    io_out_stage2Out_fixedMissPred_11=value;
  endfunction

  function void get_io_out_stage2Out_fixedMissPred_12xxPfBDHPCKVf7;
    output logic  value;
    value=io_out_stage2Out_fixedMissPred_12;
  endfunction

  function void set_io_out_stage2Out_fixedMissPred_12xxPfBDHPCKVf7;
    input logic  value;
    io_out_stage2Out_fixedMissPred_12=value;
  endfunction

  function void get_io_out_stage2Out_fixedMissPred_13xxPfBDHPCKVf7;
    output logic  value;
    value=io_out_stage2Out_fixedMissPred_13;
  endfunction

  function void set_io_out_stage2Out_fixedMissPred_13xxPfBDHPCKVf7;
    input logic  value;
    io_out_stage2Out_fixedMissPred_13=value;
  endfunction

  function void get_io_out_stage2Out_fixedMissPred_14xxPfBDHPCKVf7;
    output logic  value;
    value=io_out_stage2Out_fixedMissPred_14;
  endfunction

  function void set_io_out_stage2Out_fixedMissPred_14xxPfBDHPCKVf7;
    input logic  value;
    io_out_stage2Out_fixedMissPred_14=value;
  endfunction

  function void get_io_out_stage2Out_fixedMissPred_15xxPfBDHPCKVf7;
    output logic  value;
    value=io_out_stage2Out_fixedMissPred_15;
  endfunction

  function void set_io_out_stage2Out_fixedMissPred_15xxPfBDHPCKVf7;
    input logic  value;
    io_out_stage2Out_fixedMissPred_15=value;
  endfunction

  function void get_PredChecker_jalFaultVec_0xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.jalFaultVec_0;
  endfunction

  function void get_PredChecker_jalFaultVec_1xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.jalFaultVec_1;
  endfunction

  function void get_PredChecker_jalFaultVec_2xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.jalFaultVec_2;
  endfunction

  function void get_PredChecker_jalFaultVec_3xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.jalFaultVec_3;
  endfunction

  function void get_PredChecker_jalFaultVec_4xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.jalFaultVec_4;
  endfunction

  function void get_PredChecker_jalFaultVec_5xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.jalFaultVec_5;
  endfunction

  function void get_PredChecker_jalFaultVec_6xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.jalFaultVec_6;
  endfunction

  function void get_PredChecker_jalFaultVec_7xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.jalFaultVec_7;
  endfunction

  function void get_PredChecker_jalFaultVec_8xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.jalFaultVec_8;
  endfunction

  function void get_PredChecker_jalFaultVec_9xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.jalFaultVec_9;
  endfunction

  function void get_PredChecker_jalFaultVec_10xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.jalFaultVec_10;
  endfunction

  function void get_PredChecker_jalFaultVec_11xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.jalFaultVec_11;
  endfunction

  function void get_PredChecker_jalFaultVec_12xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.jalFaultVec_12;
  endfunction

  function void get_PredChecker_jalFaultVec_13xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.jalFaultVec_13;
  endfunction

  function void get_PredChecker_jalFaultVec_14xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.jalFaultVec_14;
  endfunction

  function void get_PredChecker_jalFaultVec_15xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.jalFaultVec_15;
  endfunction

  function void get_PredChecker_retFaultVec_0xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.retFaultVec_0;
  endfunction

  function void get_PredChecker_retFaultVec_1xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.retFaultVec_1;
  endfunction

  function void get_PredChecker_retFaultVec_2xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.retFaultVec_2;
  endfunction

  function void get_PredChecker_retFaultVec_3xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.retFaultVec_3;
  endfunction

  function void get_PredChecker_retFaultVec_4xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.retFaultVec_4;
  endfunction

  function void get_PredChecker_retFaultVec_5xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.retFaultVec_5;
  endfunction

  function void get_PredChecker_retFaultVec_6xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.retFaultVec_6;
  endfunction

  function void get_PredChecker_retFaultVec_7xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.retFaultVec_7;
  endfunction

  function void get_PredChecker_retFaultVec_8xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.retFaultVec_8;
  endfunction

  function void get_PredChecker_retFaultVec_9xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.retFaultVec_9;
  endfunction

  function void get_PredChecker_retFaultVec_10xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.retFaultVec_10;
  endfunction

  function void get_PredChecker_retFaultVec_11xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.retFaultVec_11;
  endfunction

  function void get_PredChecker_retFaultVec_12xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.retFaultVec_12;
  endfunction

  function void get_PredChecker_retFaultVec_13xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.retFaultVec_13;
  endfunction

  function void get_PredChecker_retFaultVec_14xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.retFaultVec_14;
  endfunction

  function void get_PredChecker_retFaultVec_15xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.retFaultVec_15;
  endfunction

  function void get_PredChecker_remaskFault_0xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.remaskFault_0;
  endfunction

  function void get_PredChecker_remaskFault_1xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.remaskFault_1;
  endfunction

  function void get_PredChecker_remaskFault_2xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.remaskFault_2;
  endfunction

  function void get_PredChecker_remaskFault_3xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.remaskFault_3;
  endfunction

  function void get_PredChecker_remaskFault_4xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.remaskFault_4;
  endfunction

  function void get_PredChecker_remaskFault_5xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.remaskFault_5;
  endfunction

  function void get_PredChecker_remaskFault_6xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.remaskFault_6;
  endfunction

  function void get_PredChecker_remaskFault_7xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.remaskFault_7;
  endfunction

  function void get_PredChecker_remaskFault_8xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.remaskFault_8;
  endfunction

  function void get_PredChecker_remaskFault_9xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.remaskFault_9;
  endfunction

  function void get_PredChecker_remaskFault_10xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.remaskFault_10;
  endfunction

  function void get_PredChecker_remaskFault_11xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.remaskFault_11;
  endfunction

  function void get_PredChecker_remaskFault_12xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.remaskFault_12;
  endfunction

  function void get_PredChecker_remaskFault_13xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.remaskFault_13;
  endfunction

  function void get_PredChecker_remaskFault_14xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.remaskFault_14;
  endfunction

  function void get_PredChecker_fixedRangexxPfBDHPCKVf7;
    output logic [15:0] value;
    value=PredChecker.fixedRange;
  endfunction

  function void get_PredChecker_fixedRangeNextxxPfBDHPCKVf7;
    output logic [15:0] value;
    value=PredChecker.fixedRangeNext;
  endfunction

  function void get_PredChecker_instrValidNext_0xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.instrValidNext_0;
  endfunction

  function void get_PredChecker_instrValidNext_1xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.instrValidNext_1;
  endfunction

  function void get_PredChecker_instrValidNext_2xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.instrValidNext_2;
  endfunction

  function void get_PredChecker_instrValidNext_3xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.instrValidNext_3;
  endfunction

  function void get_PredChecker_instrValidNext_4xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.instrValidNext_4;
  endfunction

  function void get_PredChecker_instrValidNext_5xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.instrValidNext_5;
  endfunction

  function void get_PredChecker_instrValidNext_6xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.instrValidNext_6;
  endfunction

  function void get_PredChecker_instrValidNext_7xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.instrValidNext_7;
  endfunction

  function void get_PredChecker_instrValidNext_8xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.instrValidNext_8;
  endfunction

  function void get_PredChecker_instrValidNext_9xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.instrValidNext_9;
  endfunction

  function void get_PredChecker_instrValidNext_10xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.instrValidNext_10;
  endfunction

  function void get_PredChecker_instrValidNext_11xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.instrValidNext_11;
  endfunction

  function void get_PredChecker_instrValidNext_12xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.instrValidNext_12;
  endfunction

  function void get_PredChecker_instrValidNext_13xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.instrValidNext_13;
  endfunction

  function void get_PredChecker_instrValidNext_14xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.instrValidNext_14;
  endfunction

  function void get_PredChecker_instrValidNext_15xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.instrValidNext_15;
  endfunction

  function void get_PredChecker_takenIdxNextxxPfBDHPCKVf7;
    output logic [3:0] value;
    value=PredChecker.takenIdxNext;
  endfunction

  function void get_PredChecker_predTakenNextxxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.predTakenNext;
  endfunction

  function void get_PredChecker_predTargetNextxxPfBDHPCKVf7;
    output logic [49:0] value;
    value=PredChecker.predTargetNext;
  endfunction

  function void get_PredChecker_jumpTargetsNext_0xxPfBDHPCKVf7;
    output logic [49:0] value;
    value=PredChecker.jumpTargetsNext_0;
  endfunction

  function void get_PredChecker_jumpTargetsNext_1xxPfBDHPCKVf7;
    output logic [49:0] value;
    value=PredChecker.jumpTargetsNext_1;
  endfunction

  function void get_PredChecker_jumpTargetsNext_2xxPfBDHPCKVf7;
    output logic [49:0] value;
    value=PredChecker.jumpTargetsNext_2;
  endfunction

  function void get_PredChecker_jumpTargetsNext_3xxPfBDHPCKVf7;
    output logic [49:0] value;
    value=PredChecker.jumpTargetsNext_3;
  endfunction

  function void get_PredChecker_jumpTargetsNext_4xxPfBDHPCKVf7;
    output logic [49:0] value;
    value=PredChecker.jumpTargetsNext_4;
  endfunction

  function void get_PredChecker_jumpTargetsNext_5xxPfBDHPCKVf7;
    output logic [49:0] value;
    value=PredChecker.jumpTargetsNext_5;
  endfunction

  function void get_PredChecker_jumpTargetsNext_6xxPfBDHPCKVf7;
    output logic [49:0] value;
    value=PredChecker.jumpTargetsNext_6;
  endfunction

  function void get_PredChecker_jumpTargetsNext_7xxPfBDHPCKVf7;
    output logic [49:0] value;
    value=PredChecker.jumpTargetsNext_7;
  endfunction

  function void get_PredChecker_jumpTargetsNext_8xxPfBDHPCKVf7;
    output logic [49:0] value;
    value=PredChecker.jumpTargetsNext_8;
  endfunction

  function void get_PredChecker_jumpTargetsNext_9xxPfBDHPCKVf7;
    output logic [49:0] value;
    value=PredChecker.jumpTargetsNext_9;
  endfunction

  function void get_PredChecker_jumpTargetsNext_10xxPfBDHPCKVf7;
    output logic [49:0] value;
    value=PredChecker.jumpTargetsNext_10;
  endfunction

  function void get_PredChecker_jumpTargetsNext_11xxPfBDHPCKVf7;
    output logic [49:0] value;
    value=PredChecker.jumpTargetsNext_11;
  endfunction

  function void get_PredChecker_jumpTargetsNext_12xxPfBDHPCKVf7;
    output logic [49:0] value;
    value=PredChecker.jumpTargetsNext_12;
  endfunction

  function void get_PredChecker_jumpTargetsNext_13xxPfBDHPCKVf7;
    output logic [49:0] value;
    value=PredChecker.jumpTargetsNext_13;
  endfunction

  function void get_PredChecker_jumpTargetsNext_14xxPfBDHPCKVf7;
    output logic [49:0] value;
    value=PredChecker.jumpTargetsNext_14;
  endfunction

  function void get_PredChecker_jumpTargetsNext_15xxPfBDHPCKVf7;
    output logic [49:0] value;
    value=PredChecker.jumpTargetsNext_15;
  endfunction

  function void get_PredChecker_seqTargetsNext_0xxPfBDHPCKVf7;
    output logic [49:0] value;
    value=PredChecker.seqTargetsNext_0;
  endfunction

  function void get_PredChecker_seqTargetsNext_1xxPfBDHPCKVf7;
    output logic [49:0] value;
    value=PredChecker.seqTargetsNext_1;
  endfunction

  function void get_PredChecker_seqTargetsNext_2xxPfBDHPCKVf7;
    output logic [49:0] value;
    value=PredChecker.seqTargetsNext_2;
  endfunction

  function void get_PredChecker_seqTargetsNext_3xxPfBDHPCKVf7;
    output logic [49:0] value;
    value=PredChecker.seqTargetsNext_3;
  endfunction

  function void get_PredChecker_seqTargetsNext_4xxPfBDHPCKVf7;
    output logic [49:0] value;
    value=PredChecker.seqTargetsNext_4;
  endfunction

  function void get_PredChecker_seqTargetsNext_5xxPfBDHPCKVf7;
    output logic [49:0] value;
    value=PredChecker.seqTargetsNext_5;
  endfunction

  function void get_PredChecker_seqTargetsNext_6xxPfBDHPCKVf7;
    output logic [49:0] value;
    value=PredChecker.seqTargetsNext_6;
  endfunction

  function void get_PredChecker_seqTargetsNext_7xxPfBDHPCKVf7;
    output logic [49:0] value;
    value=PredChecker.seqTargetsNext_7;
  endfunction

  function void get_PredChecker_seqTargetsNext_8xxPfBDHPCKVf7;
    output logic [49:0] value;
    value=PredChecker.seqTargetsNext_8;
  endfunction

  function void get_PredChecker_seqTargetsNext_9xxPfBDHPCKVf7;
    output logic [49:0] value;
    value=PredChecker.seqTargetsNext_9;
  endfunction

  function void get_PredChecker_seqTargetsNext_10xxPfBDHPCKVf7;
    output logic [49:0] value;
    value=PredChecker.seqTargetsNext_10;
  endfunction

  function void get_PredChecker_seqTargetsNext_11xxPfBDHPCKVf7;
    output logic [49:0] value;
    value=PredChecker.seqTargetsNext_11;
  endfunction

  function void get_PredChecker_seqTargetsNext_12xxPfBDHPCKVf7;
    output logic [49:0] value;
    value=PredChecker.seqTargetsNext_12;
  endfunction

  function void get_PredChecker_seqTargetsNext_13xxPfBDHPCKVf7;
    output logic [49:0] value;
    value=PredChecker.seqTargetsNext_13;
  endfunction

  function void get_PredChecker_seqTargetsNext_14xxPfBDHPCKVf7;
    output logic [49:0] value;
    value=PredChecker.seqTargetsNext_14;
  endfunction

  function void get_PredChecker_seqTargetsNext_15xxPfBDHPCKVf7;
    output logic [49:0] value;
    value=PredChecker.seqTargetsNext_15;
  endfunction

  function void get_PredChecker_pdsNext_0_brTypexxPfBDHPCKVf7;
    output logic [1:0] value;
    value=PredChecker.pdsNext_0_brType;
  endfunction

  function void get_PredChecker_pdsNext_1_brTypexxPfBDHPCKVf7;
    output logic [1:0] value;
    value=PredChecker.pdsNext_1_brType;
  endfunction

  function void get_PredChecker_pdsNext_2_brTypexxPfBDHPCKVf7;
    output logic [1:0] value;
    value=PredChecker.pdsNext_2_brType;
  endfunction

  function void get_PredChecker_pdsNext_3_brTypexxPfBDHPCKVf7;
    output logic [1:0] value;
    value=PredChecker.pdsNext_3_brType;
  endfunction

  function void get_PredChecker_pdsNext_4_brTypexxPfBDHPCKVf7;
    output logic [1:0] value;
    value=PredChecker.pdsNext_4_brType;
  endfunction

  function void get_PredChecker_pdsNext_5_brTypexxPfBDHPCKVf7;
    output logic [1:0] value;
    value=PredChecker.pdsNext_5_brType;
  endfunction

  function void get_PredChecker_pdsNext_6_brTypexxPfBDHPCKVf7;
    output logic [1:0] value;
    value=PredChecker.pdsNext_6_brType;
  endfunction

  function void get_PredChecker_pdsNext_7_brTypexxPfBDHPCKVf7;
    output logic [1:0] value;
    value=PredChecker.pdsNext_7_brType;
  endfunction

  function void get_PredChecker_pdsNext_8_brTypexxPfBDHPCKVf7;
    output logic [1:0] value;
    value=PredChecker.pdsNext_8_brType;
  endfunction

  function void get_PredChecker_pdsNext_9_brTypexxPfBDHPCKVf7;
    output logic [1:0] value;
    value=PredChecker.pdsNext_9_brType;
  endfunction

  function void get_PredChecker_pdsNext_10_brTypexxPfBDHPCKVf7;
    output logic [1:0] value;
    value=PredChecker.pdsNext_10_brType;
  endfunction

  function void get_PredChecker_pdsNext_11_brTypexxPfBDHPCKVf7;
    output logic [1:0] value;
    value=PredChecker.pdsNext_11_brType;
  endfunction

  function void get_PredChecker_pdsNext_12_brTypexxPfBDHPCKVf7;
    output logic [1:0] value;
    value=PredChecker.pdsNext_12_brType;
  endfunction

  function void get_PredChecker_pdsNext_13_brTypexxPfBDHPCKVf7;
    output logic [1:0] value;
    value=PredChecker.pdsNext_13_brType;
  endfunction

  function void get_PredChecker_pdsNext_14_brTypexxPfBDHPCKVf7;
    output logic [1:0] value;
    value=PredChecker.pdsNext_14_brType;
  endfunction

  function void get_PredChecker_pdsNext_15_brTypexxPfBDHPCKVf7;
    output logic [1:0] value;
    value=PredChecker.pdsNext_15_brType;
  endfunction

  function void get_PredChecker_jalFaultVecNext_0xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.jalFaultVecNext_0;
  endfunction

  function void get_PredChecker_jalFaultVecNext_1xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.jalFaultVecNext_1;
  endfunction

  function void get_PredChecker_jalFaultVecNext_2xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.jalFaultVecNext_2;
  endfunction

  function void get_PredChecker_jalFaultVecNext_3xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.jalFaultVecNext_3;
  endfunction

  function void get_PredChecker_jalFaultVecNext_4xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.jalFaultVecNext_4;
  endfunction

  function void get_PredChecker_jalFaultVecNext_5xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.jalFaultVecNext_5;
  endfunction

  function void get_PredChecker_jalFaultVecNext_6xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.jalFaultVecNext_6;
  endfunction

  function void get_PredChecker_jalFaultVecNext_7xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.jalFaultVecNext_7;
  endfunction

  function void get_PredChecker_jalFaultVecNext_8xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.jalFaultVecNext_8;
  endfunction

  function void get_PredChecker_jalFaultVecNext_9xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.jalFaultVecNext_9;
  endfunction

  function void get_PredChecker_jalFaultVecNext_10xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.jalFaultVecNext_10;
  endfunction

  function void get_PredChecker_jalFaultVecNext_11xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.jalFaultVecNext_11;
  endfunction

  function void get_PredChecker_jalFaultVecNext_12xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.jalFaultVecNext_12;
  endfunction

  function void get_PredChecker_jalFaultVecNext_13xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.jalFaultVecNext_13;
  endfunction

  function void get_PredChecker_jalFaultVecNext_14xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.jalFaultVecNext_14;
  endfunction

  function void get_PredChecker_jalFaultVecNext_15xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.jalFaultVecNext_15;
  endfunction

  function void get_PredChecker_retFaultVecNext_0xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.retFaultVecNext_0;
  endfunction

  function void get_PredChecker_retFaultVecNext_1xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.retFaultVecNext_1;
  endfunction

  function void get_PredChecker_retFaultVecNext_2xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.retFaultVecNext_2;
  endfunction

  function void get_PredChecker_retFaultVecNext_3xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.retFaultVecNext_3;
  endfunction

  function void get_PredChecker_retFaultVecNext_4xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.retFaultVecNext_4;
  endfunction

  function void get_PredChecker_retFaultVecNext_5xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.retFaultVecNext_5;
  endfunction

  function void get_PredChecker_retFaultVecNext_6xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.retFaultVecNext_6;
  endfunction

  function void get_PredChecker_retFaultVecNext_7xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.retFaultVecNext_7;
  endfunction

  function void get_PredChecker_retFaultVecNext_8xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.retFaultVecNext_8;
  endfunction

  function void get_PredChecker_retFaultVecNext_9xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.retFaultVecNext_9;
  endfunction

  function void get_PredChecker_retFaultVecNext_10xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.retFaultVecNext_10;
  endfunction

  function void get_PredChecker_retFaultVecNext_11xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.retFaultVecNext_11;
  endfunction

  function void get_PredChecker_retFaultVecNext_12xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.retFaultVecNext_12;
  endfunction

  function void get_PredChecker_retFaultVecNext_13xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.retFaultVecNext_13;
  endfunction

  function void get_PredChecker_retFaultVecNext_14xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.retFaultVecNext_14;
  endfunction

  function void get_PredChecker_retFaultVecNext_15xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.retFaultVecNext_15;
  endfunction

  function void get_PredChecker_notCFITakenNext_0xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.notCFITakenNext_0;
  endfunction

  function void get_PredChecker_notCFITakenNext_1xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.notCFITakenNext_1;
  endfunction

  function void get_PredChecker_notCFITakenNext_2xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.notCFITakenNext_2;
  endfunction

  function void get_PredChecker_notCFITakenNext_3xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.notCFITakenNext_3;
  endfunction

  function void get_PredChecker_notCFITakenNext_4xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.notCFITakenNext_4;
  endfunction

  function void get_PredChecker_notCFITakenNext_5xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.notCFITakenNext_5;
  endfunction

  function void get_PredChecker_notCFITakenNext_6xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.notCFITakenNext_6;
  endfunction

  function void get_PredChecker_notCFITakenNext_7xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.notCFITakenNext_7;
  endfunction

  function void get_PredChecker_notCFITakenNext_8xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.notCFITakenNext_8;
  endfunction

  function void get_PredChecker_notCFITakenNext_9xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.notCFITakenNext_9;
  endfunction

  function void get_PredChecker_notCFITakenNext_10xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.notCFITakenNext_10;
  endfunction

  function void get_PredChecker_notCFITakenNext_11xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.notCFITakenNext_11;
  endfunction

  function void get_PredChecker_notCFITakenNext_12xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.notCFITakenNext_12;
  endfunction

  function void get_PredChecker_notCFITakenNext_13xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.notCFITakenNext_13;
  endfunction

  function void get_PredChecker_notCFITakenNext_14xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.notCFITakenNext_14;
  endfunction

  function void get_PredChecker_notCFITakenNext_15xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.notCFITakenNext_15;
  endfunction

  function void get_PredChecker_invalidTakenNext_0xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.invalidTakenNext_0;
  endfunction

  function void get_PredChecker_invalidTakenNext_1xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.invalidTakenNext_1;
  endfunction

  function void get_PredChecker_invalidTakenNext_2xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.invalidTakenNext_2;
  endfunction

  function void get_PredChecker_invalidTakenNext_3xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.invalidTakenNext_3;
  endfunction

  function void get_PredChecker_invalidTakenNext_4xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.invalidTakenNext_4;
  endfunction

  function void get_PredChecker_invalidTakenNext_5xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.invalidTakenNext_5;
  endfunction

  function void get_PredChecker_invalidTakenNext_6xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.invalidTakenNext_6;
  endfunction

  function void get_PredChecker_invalidTakenNext_7xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.invalidTakenNext_7;
  endfunction

  function void get_PredChecker_invalidTakenNext_8xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.invalidTakenNext_8;
  endfunction

  function void get_PredChecker_invalidTakenNext_9xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.invalidTakenNext_9;
  endfunction

  function void get_PredChecker_invalidTakenNext_10xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.invalidTakenNext_10;
  endfunction

  function void get_PredChecker_invalidTakenNext_11xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.invalidTakenNext_11;
  endfunction

  function void get_PredChecker_invalidTakenNext_12xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.invalidTakenNext_12;
  endfunction

  function void get_PredChecker_invalidTakenNext_13xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.invalidTakenNext_13;
  endfunction

  function void get_PredChecker_invalidTakenNext_14xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.invalidTakenNext_14;
  endfunction

  function void get_PredChecker_invalidTakenNext_15xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.invalidTakenNext_15;
  endfunction

  function void get_PredChecker_targetFault_0xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.targetFault_0;
  endfunction

  function void get_PredChecker_targetFault_1xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.targetFault_1;
  endfunction

  function void get_PredChecker_targetFault_2xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.targetFault_2;
  endfunction

  function void get_PredChecker_targetFault_3xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.targetFault_3;
  endfunction

  function void get_PredChecker_targetFault_4xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.targetFault_4;
  endfunction

  function void get_PredChecker_targetFault_5xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.targetFault_5;
  endfunction

  function void get_PredChecker_targetFault_6xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.targetFault_6;
  endfunction

  function void get_PredChecker_targetFault_7xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.targetFault_7;
  endfunction

  function void get_PredChecker_targetFault_8xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.targetFault_8;
  endfunction

  function void get_PredChecker_targetFault_9xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.targetFault_9;
  endfunction

  function void get_PredChecker_targetFault_10xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.targetFault_10;
  endfunction

  function void get_PredChecker_targetFault_11xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.targetFault_11;
  endfunction

  function void get_PredChecker_targetFault_12xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.targetFault_12;
  endfunction

  function void get_PredChecker_targetFault_13xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.targetFault_13;
  endfunction

  function void get_PredChecker_targetFault_14xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.targetFault_14;
  endfunction

  function void get_PredChecker_targetFault_15xxPfBDHPCKVf7;
    output logic  value;
    value=PredChecker.targetFault_15;
  endfunction



  initial begin
    $dumpfile("PredChecker.fst");
    $dumpvars(0, PredChecker_top);
  end

  export "DPI-C" function finish_PfBDHPCKVf7;
  function void finish_PfBDHPCKVf7;
    $finish;
  endfunction


endmodule
